module system_top (ref_clk, uart_clk, reset_n, rx_in, tx_out);

input ref_clk;
input uart_clk;
input reset_n;
input rx_in;
output tx_out;

wire vdd = 1'b1;
wire gnd = 1'b0;

INVX1 INVX1_1 ( .A(alu_inst_alu_out_comp_valid), .Y(_406_) );
INVX1 INVX1_2 ( .A(alu_inst_alu_func_in_1_), .Y(_417_) );
INVX1 INVX1_3 ( .A(alu_inst_alu_func_in_0_), .Y(_428_) );
NOR2X1 NOR2X1_1 ( .A(_417_), .B(_428_), .Y(_439_) );
INVX1 INVX1_4 ( .A(_439_), .Y(_450_) );
NOR2X1 NOR2X1_2 ( .A(alu_inst_alu_func_in_2_), .B(alu_inst_alu_func_in_3_), .Y(_461_) );
INVX1 INVX1_5 ( .A(_461_), .Y(_472_) );
NOR2X1 NOR2X1_3 ( .A(_472_), .B(_450_), .Y(_483_) );
NOR2X1 NOR2X1_4 ( .A(alu_inst_data_b_in_4_), .B(alu_inst_data_b_in_3_), .Y(_494_) );
INVX1 INVX1_6 ( .A(alu_inst_data_b_in_5_), .Y(_505_) );
NOR2X1 NOR2X1_5 ( .A(alu_inst_data_b_in_7_), .B(alu_inst_data_b_in_6_), .Y(_516_) );
AND2X2 AND2X2_1 ( .A(_516_), .B(_505_), .Y(_527_) );
NAND2X1 NAND2X1_1 ( .A(_494_), .B(_527_), .Y(_538_) );
INVX1 INVX1_7 ( .A(alu_inst_data_b_in_2_), .Y(_549_) );
INVX1 INVX1_8 ( .A(alu_inst_data_a_in_7_), .Y(_560_) );
INVX1 INVX1_9 ( .A(alu_inst_data_b_in_0_), .Y(_571_) );
INVX1 INVX1_10 ( .A(alu_inst_data_b_in_7_), .Y(_582_) );
INVX1 INVX1_11 ( .A(alu_inst_data_b_in_6_), .Y(_593_) );
NAND3X1 NAND3X1_1 ( .A(_582_), .B(_593_), .C(_505_), .Y(_604_) );
NOR2X1 NOR2X1_6 ( .A(alu_inst_data_b_in_2_), .B(alu_inst_data_b_in_1_), .Y(_614_) );
NAND2X1 NAND2X1_2 ( .A(_494_), .B(_614_), .Y(_625_) );
NOR3X1 NOR3X1_1 ( .A(_571_), .B(_604_), .C(_625_), .Y(_636_) );
NOR2X1 NOR2X1_7 ( .A(_560_), .B(_636_), .Y(_646_) );
NAND3X1 NAND3X1_2 ( .A(_549_), .B(_494_), .C(_527_), .Y(_657_) );
INVX1 INVX1_12 ( .A(_657_), .Y(_668_) );
INVX1 INVX1_13 ( .A(alu_inst_data_b_in_1_), .Y(_679_) );
OAI21X1 OAI21X1_1 ( .A(alu_inst_data_a_in_6_), .B(_571_), .C(_679_), .Y(_689_) );
NOR2X1 NOR2X1_8 ( .A(alu_inst_data_a_in_6_), .B(_571_), .Y(_700_) );
NAND2X1 NAND2X1_3 ( .A(alu_inst_data_b_in_1_), .B(_700_), .Y(_711_) );
NAND3X1 NAND3X1_3 ( .A(_689_), .B(_711_), .C(_668_), .Y(_721_) );
NAND3X1 NAND3X1_4 ( .A(_549_), .B(_646_), .C(_721_), .Y(_732_) );
OAI21X1 OAI21X1_2 ( .A(_549_), .B(_646_), .C(_732_), .Y(_743_) );
INVX1 INVX1_14 ( .A(_743_), .Y(_754_) );
OAI21X1 OAI21X1_3 ( .A(_560_), .B(_636_), .C(_689_), .Y(_765_) );
AOI21X1 AOI21X1_1 ( .A(alu_inst_data_b_in_1_), .B(_700_), .C(_657_), .Y(_775_) );
NAND3X1 NAND3X1_5 ( .A(alu_inst_data_b_in_0_), .B(_775_), .C(_765_), .Y(_786_) );
NAND3X1 NAND3X1_6 ( .A(alu_inst_data_a_in_6_), .B(_679_), .C(_786_), .Y(_797_) );
AOI21X1 AOI21X1_2 ( .A(_786_), .B(alu_inst_data_a_in_6_), .C(_679_), .Y(_808_) );
INVX1 INVX1_15 ( .A(alu_inst_data_a_in_5_), .Y(_818_) );
NOR2X1 NOR2X1_9 ( .A(alu_inst_data_a_in_4_), .B(_571_), .Y(_829_) );
INVX1 INVX1_16 ( .A(alu_inst_data_a_in_4_), .Y(_840_) );
NOR2X1 NOR2X1_10 ( .A(_840_), .B(_571_), .Y(_851_) );
INVX1 INVX1_17 ( .A(_851_), .Y(_862_) );
XNOR2X1 XNOR2X1_1 ( .A(alu_inst_data_a_in_5_), .B(alu_inst_data_b_in_0_), .Y(_873_) );
OAI21X1 OAI21X1_4 ( .A(alu_inst_data_a_in_4_), .B(_873_), .C(_862_), .Y(_884_) );
OAI21X1 OAI21X1_5 ( .A(_818_), .B(_829_), .C(_884_), .Y(_894_) );
INVX1 INVX1_18 ( .A(_894_), .Y(_905_) );
OAI21X1 OAI21X1_6 ( .A(_905_), .B(_808_), .C(_797_), .Y(_916_) );
NAND2X1 NAND2X1_4 ( .A(_754_), .B(_916_), .Y(_927_) );
AOI21X1 AOI21X1_3 ( .A(_927_), .B(_732_), .C(_538_), .Y(_938_) );
XNOR2X1 XNOR2X1_2 ( .A(_916_), .B(_743_), .Y(_949_) );
NAND2X1 NAND2X1_5 ( .A(_949_), .B(_938_), .Y(_959_) );
INVX1 INVX1_19 ( .A(_959_), .Y(_970_) );
INVX1 INVX1_20 ( .A(_538_), .Y(_981_) );
NAND2X1 NAND2X1_6 ( .A(_732_), .B(_927_), .Y(_992_) );
NAND2X1 NAND2X1_7 ( .A(_981_), .B(_992_), .Y(_1003_) );
NAND2X1 NAND2X1_8 ( .A(_646_), .B(_721_), .Y(_1014_) );
INVX1 INVX1_21 ( .A(_732_), .Y(_1024_) );
AOI21X1 AOI21X1_4 ( .A(_916_), .B(_754_), .C(_1024_), .Y(_1035_) );
OAI21X1 OAI21X1_7 ( .A(_538_), .B(_1035_), .C(_1014_), .Y(_1046_) );
OAI21X1 OAI21X1_8 ( .A(_949_), .B(_1003_), .C(_1046_), .Y(_1057_) );
NOR2X1 NOR2X1_11 ( .A(alu_inst_data_b_in_4_), .B(_604_), .Y(_1067_) );
NAND2X1 NAND2X1_9 ( .A(alu_inst_data_a_in_6_), .B(_786_), .Y(_10_) );
NAND2X1 NAND2X1_10 ( .A(alu_inst_data_b_in_1_), .B(_10_), .Y(_21_) );
NAND3X1 NAND3X1_7 ( .A(_797_), .B(_894_), .C(_21_), .Y(_32_) );
INVX1 INVX1_22 ( .A(_797_), .Y(_42_) );
OAI21X1 OAI21X1_9 ( .A(_808_), .B(_42_), .C(_905_), .Y(_53_) );
NAND2X1 NAND2X1_11 ( .A(_32_), .B(_53_), .Y(_63_) );
NAND3X1 NAND3X1_8 ( .A(_981_), .B(_63_), .C(_992_), .Y(_74_) );
OAI21X1 OAI21X1_10 ( .A(_538_), .B(_1035_), .C(_10_), .Y(_85_) );
NAND3X1 NAND3X1_9 ( .A(_549_), .B(_85_), .C(_74_), .Y(_95_) );
INVX1 INVX1_23 ( .A(_95_), .Y(_106_) );
XOR2X1 XOR2X1_1 ( .A(_916_), .B(_743_), .Y(_116_) );
NAND2X1 NAND2X1_12 ( .A(_116_), .B(_938_), .Y(_126_) );
NAND3X1 NAND3X1_10 ( .A(alu_inst_data_b_in_3_), .B(_1046_), .C(_126_), .Y(_128_) );
INVX1 INVX1_24 ( .A(alu_inst_data_b_in_3_), .Y(_129_) );
INVX1 INVX1_25 ( .A(_1014_), .Y(_130_) );
OAI21X1 OAI21X1_11 ( .A(_538_), .B(_1035_), .C(_130_), .Y(_131_) );
NAND3X1 NAND3X1_11 ( .A(_129_), .B(_131_), .C(_959_), .Y(_132_) );
NAND2X1 NAND2X1_13 ( .A(_128_), .B(_132_), .Y(_133_) );
AOI21X1 AOI21X1_5 ( .A(_959_), .B(_131_), .C(alu_inst_data_b_in_3_), .Y(_134_) );
AOI21X1 AOI21X1_6 ( .A(_133_), .B(_106_), .C(_134_), .Y(_135_) );
AND2X2 AND2X2_2 ( .A(_53_), .B(_32_), .Y(_136_) );
NAND3X1 NAND3X1_12 ( .A(_981_), .B(_992_), .C(_136_), .Y(_137_) );
INVX1 INVX1_26 ( .A(_10_), .Y(_138_) );
OAI21X1 OAI21X1_12 ( .A(_538_), .B(_1035_), .C(_138_), .Y(_139_) );
NAND3X1 NAND3X1_13 ( .A(alu_inst_data_b_in_2_), .B(_139_), .C(_137_), .Y(_140_) );
AND2X2 AND2X2_3 ( .A(_140_), .B(_95_), .Y(_141_) );
NAND3X1 NAND3X1_14 ( .A(_981_), .B(_873_), .C(_992_), .Y(_142_) );
OAI21X1 OAI21X1_13 ( .A(_538_), .B(_1035_), .C(_818_), .Y(_143_) );
NAND3X1 NAND3X1_15 ( .A(_679_), .B(_143_), .C(_142_), .Y(_144_) );
AOI21X1 AOI21X1_7 ( .A(_142_), .B(_143_), .C(_679_), .Y(_145_) );
OAI21X1 OAI21X1_14 ( .A(_829_), .B(_145_), .C(_144_), .Y(_146_) );
NAND3X1 NAND3X1_16 ( .A(_133_), .B(_141_), .C(_146_), .Y(_147_) );
NAND2X1 NAND2X1_14 ( .A(_135_), .B(_147_), .Y(_148_) );
AOI21X1 AOI21X1_8 ( .A(_148_), .B(_1067_), .C(_1057_), .Y(_149_) );
NOR2X1 NOR2X1_12 ( .A(_970_), .B(_149_), .Y(_150_) );
INVX1 INVX1_27 ( .A(_150_), .Y(_151_) );
INVX1 INVX1_28 ( .A(alu_inst_data_b_in_4_), .Y(_152_) );
XNOR2X1 XNOR2X1_3 ( .A(_146_), .B(_141_), .Y(_153_) );
NAND3X1 NAND3X1_17 ( .A(_1067_), .B(_148_), .C(_153_), .Y(_154_) );
INVX1 INVX1_29 ( .A(_1067_), .Y(_155_) );
OAI21X1 OAI21X1_15 ( .A(_138_), .B(_938_), .C(_74_), .Y(_156_) );
AND2X2 AND2X2_4 ( .A(_147_), .B(_135_), .Y(_157_) );
OAI21X1 OAI21X1_16 ( .A(_155_), .B(_157_), .C(_156_), .Y(_158_) );
NAND3X1 NAND3X1_18 ( .A(_129_), .B(_154_), .C(_158_), .Y(_159_) );
OAI21X1 OAI21X1_17 ( .A(alu_inst_data_b_in_4_), .B(_150_), .C(_159_), .Y(_160_) );
OAI21X1 OAI21X1_18 ( .A(_152_), .B(_151_), .C(_160_), .Y(_161_) );
OAI21X1 OAI21X1_19 ( .A(_970_), .B(_149_), .C(alu_inst_data_b_in_4_), .Y(_162_) );
NAND2X1 NAND2X1_15 ( .A(_152_), .B(_150_), .Y(_163_) );
XOR2X1 XOR2X1_2 ( .A(_146_), .B(_141_), .Y(_164_) );
NAND3X1 NAND3X1_19 ( .A(_1067_), .B(_148_), .C(_164_), .Y(_165_) );
INVX1 INVX1_30 ( .A(_156_), .Y(_166_) );
OAI21X1 OAI21X1_20 ( .A(_155_), .B(_157_), .C(_166_), .Y(_167_) );
NAND3X1 NAND3X1_20 ( .A(alu_inst_data_b_in_3_), .B(_165_), .C(_167_), .Y(_168_) );
NAND2X1 NAND2X1_16 ( .A(_159_), .B(_168_), .Y(_169_) );
AOI21X1 AOI21X1_9 ( .A(_162_), .B(_163_), .C(_169_), .Y(_170_) );
AND2X2 AND2X2_5 ( .A(_142_), .B(_143_), .Y(_171_) );
OAI21X1 OAI21X1_21 ( .A(_155_), .B(_157_), .C(_171_), .Y(_172_) );
NAND2X1 NAND2X1_17 ( .A(alu_inst_data_b_in_1_), .B(_171_), .Y(_173_) );
OAI21X1 OAI21X1_22 ( .A(alu_inst_data_a_in_5_), .B(_938_), .C(_142_), .Y(_174_) );
NAND2X1 NAND2X1_18 ( .A(_679_), .B(_174_), .Y(_175_) );
NAND2X1 NAND2X1_19 ( .A(_175_), .B(_173_), .Y(_176_) );
OAI21X1 OAI21X1_23 ( .A(alu_inst_data_a_in_4_), .B(_571_), .C(_176_), .Y(_177_) );
NAND3X1 NAND3X1_21 ( .A(_829_), .B(_175_), .C(_173_), .Y(_178_) );
AND2X2 AND2X2_6 ( .A(_177_), .B(_178_), .Y(_179_) );
NAND3X1 NAND3X1_22 ( .A(_1067_), .B(_148_), .C(_179_), .Y(_180_) );
NAND3X1 NAND3X1_23 ( .A(alu_inst_data_b_in_2_), .B(_172_), .C(_180_), .Y(_181_) );
NAND2X1 NAND2X1_20 ( .A(_1067_), .B(_148_), .Y(_182_) );
NAND2X1 NAND2X1_21 ( .A(_178_), .B(_177_), .Y(_183_) );
OAI21X1 OAI21X1_24 ( .A(_182_), .B(_183_), .C(_172_), .Y(_184_) );
NAND2X1 NAND2X1_22 ( .A(_549_), .B(_184_), .Y(_185_) );
NOR2X1 NOR2X1_13 ( .A(alu_inst_data_b_in_0_), .B(_840_), .Y(_186_) );
NOR2X1 NOR2X1_14 ( .A(_829_), .B(_186_), .Y(_187_) );
NAND3X1 NAND3X1_24 ( .A(_1067_), .B(_187_), .C(_148_), .Y(_188_) );
OAI21X1 OAI21X1_25 ( .A(_155_), .B(_157_), .C(_840_), .Y(_189_) );
NAND3X1 NAND3X1_25 ( .A(_679_), .B(_188_), .C(_189_), .Y(_190_) );
NOR2X1 NOR2X1_15 ( .A(alu_inst_data_a_in_3_), .B(_571_), .Y(_191_) );
INVX1 INVX1_31 ( .A(_191_), .Y(_192_) );
NAND2X1 NAND2X1_23 ( .A(alu_inst_data_b_in_0_), .B(_1067_), .Y(_193_) );
OAI21X1 OAI21X1_26 ( .A(_193_), .B(_157_), .C(alu_inst_data_a_in_4_), .Y(_194_) );
INVX1 INVX1_32 ( .A(_193_), .Y(_195_) );
NAND3X1 NAND3X1_26 ( .A(_840_), .B(_195_), .C(_148_), .Y(_196_) );
NAND3X1 NAND3X1_27 ( .A(alu_inst_data_b_in_1_), .B(_196_), .C(_194_), .Y(_197_) );
NAND3X1 NAND3X1_28 ( .A(_192_), .B(_190_), .C(_197_), .Y(_198_) );
NAND3X1 NAND3X1_29 ( .A(_185_), .B(_190_), .C(_198_), .Y(_199_) );
NAND3X1 NAND3X1_30 ( .A(_181_), .B(_199_), .C(_170_), .Y(_200_) );
AOI21X1 AOI21X1_10 ( .A(_200_), .B(_161_), .C(_604_), .Y(_201_) );
NAND2X1 NAND2X1_24 ( .A(_162_), .B(_163_), .Y(_202_) );
INVX1 INVX1_33 ( .A(_169_), .Y(_203_) );
INVX1 INVX1_34 ( .A(_181_), .Y(_204_) );
AOI21X1 AOI21X1_11 ( .A(_194_), .B(_196_), .C(alu_inst_data_b_in_1_), .Y(_205_) );
AOI21X1 AOI21X1_12 ( .A(_192_), .B(_197_), .C(_205_), .Y(_206_) );
OAI21X1 OAI21X1_27 ( .A(_204_), .B(_206_), .C(_185_), .Y(_207_) );
NAND2X1 NAND2X1_25 ( .A(_203_), .B(_207_), .Y(_208_) );
NAND3X1 NAND3X1_31 ( .A(_159_), .B(_202_), .C(_208_), .Y(_209_) );
INVX1 INVX1_35 ( .A(_159_), .Y(_210_) );
INVX1 INVX1_36 ( .A(_202_), .Y(_211_) );
AOI21X1 AOI21X1_13 ( .A(_180_), .B(_172_), .C(alu_inst_data_b_in_2_), .Y(_212_) );
AOI21X1 AOI21X1_14 ( .A(_181_), .B(_205_), .C(_212_), .Y(_213_) );
AND2X2 AND2X2_7 ( .A(_190_), .B(_197_), .Y(_214_) );
NAND3X1 NAND3X1_32 ( .A(_1067_), .B(_148_), .C(_183_), .Y(_215_) );
OAI21X1 OAI21X1_28 ( .A(_155_), .B(_157_), .C(_174_), .Y(_216_) );
NAND3X1 NAND3X1_33 ( .A(alu_inst_data_b_in_2_), .B(_215_), .C(_216_), .Y(_217_) );
NAND3X1 NAND3X1_34 ( .A(_549_), .B(_172_), .C(_180_), .Y(_218_) );
NAND2X1 NAND2X1_26 ( .A(_217_), .B(_218_), .Y(_219_) );
NAND3X1 NAND3X1_35 ( .A(_192_), .B(_219_), .C(_214_), .Y(_220_) );
AOI21X1 AOI21X1_15 ( .A(_220_), .B(_213_), .C(_169_), .Y(_221_) );
OAI21X1 OAI21X1_29 ( .A(_210_), .B(_221_), .C(_211_), .Y(_222_) );
NAND3X1 NAND3X1_36 ( .A(_201_), .B(_209_), .C(_222_), .Y(_223_) );
OAI21X1 OAI21X1_30 ( .A(_151_), .B(_201_), .C(_223_), .Y(_224_) );
INVX1 INVX1_37 ( .A(_516_), .Y(_225_) );
NAND2X1 NAND2X1_27 ( .A(alu_inst_data_b_in_4_), .B(_150_), .Y(_226_) );
AOI22X1 AOI22X1_1 ( .A(_226_), .B(_160_), .C(_207_), .D(_170_), .Y(_227_) );
OAI21X1 OAI21X1_31 ( .A(_604_), .B(_227_), .C(_150_), .Y(_228_) );
NAND3X1 NAND3X1_37 ( .A(_505_), .B(_228_), .C(_223_), .Y(_229_) );
NOR2X1 NOR2X1_16 ( .A(_203_), .B(_207_), .Y(_230_) );
OAI21X1 OAI21X1_32 ( .A(_221_), .B(_230_), .C(_201_), .Y(_231_) );
OAI21X1 OAI21X1_33 ( .A(_182_), .B(_164_), .C(_158_), .Y(_232_) );
OAI21X1 OAI21X1_34 ( .A(_604_), .B(_227_), .C(_232_), .Y(_233_) );
NAND3X1 NAND3X1_38 ( .A(_152_), .B(_233_), .C(_231_), .Y(_234_) );
AOI21X1 AOI21X1_16 ( .A(_223_), .B(_228_), .C(_505_), .Y(_235_) );
OAI21X1 OAI21X1_35 ( .A(_234_), .B(_235_), .C(_229_), .Y(_236_) );
NAND3X1 NAND3X1_39 ( .A(alu_inst_data_b_in_5_), .B(_228_), .C(_223_), .Y(_237_) );
INVX1 INVX1_38 ( .A(_228_), .Y(_238_) );
NAND2X1 NAND2X1_28 ( .A(_202_), .B(_203_), .Y(_239_) );
AOI21X1 AOI21X1_17 ( .A(_189_), .B(_188_), .C(_679_), .Y(_240_) );
OAI21X1 OAI21X1_36 ( .A(_191_), .B(_240_), .C(_190_), .Y(_241_) );
AOI21X1 AOI21X1_18 ( .A(_241_), .B(_181_), .C(_212_), .Y(_242_) );
OAI21X1 OAI21X1_37 ( .A(_239_), .B(_242_), .C(_161_), .Y(_243_) );
NAND2X1 NAND2X1_29 ( .A(_527_), .B(_243_), .Y(_244_) );
NAND3X1 NAND3X1_40 ( .A(_159_), .B(_211_), .C(_208_), .Y(_245_) );
OAI21X1 OAI21X1_38 ( .A(_210_), .B(_221_), .C(_202_), .Y(_246_) );
AOI21X1 AOI21X1_19 ( .A(_246_), .B(_245_), .C(_244_), .Y(_247_) );
OAI21X1 OAI21X1_39 ( .A(_238_), .B(_247_), .C(_505_), .Y(_248_) );
NAND2X1 NAND2X1_30 ( .A(_169_), .B(_242_), .Y(_249_) );
NAND3X1 NAND3X1_41 ( .A(_208_), .B(_249_), .C(_201_), .Y(_250_) );
INVX1 INVX1_39 ( .A(_232_), .Y(_251_) );
OAI21X1 OAI21X1_40 ( .A(_604_), .B(_227_), .C(_251_), .Y(_252_) );
NAND3X1 NAND3X1_42 ( .A(alu_inst_data_b_in_4_), .B(_252_), .C(_250_), .Y(_253_) );
NAND2X1 NAND2X1_31 ( .A(_234_), .B(_253_), .Y(_254_) );
AOI21X1 AOI21X1_20 ( .A(_237_), .B(_248_), .C(_254_), .Y(_255_) );
XNOR2X1 XNOR2X1_4 ( .A(_241_), .B(_219_), .Y(_256_) );
NAND3X1 NAND3X1_43 ( .A(_527_), .B(_256_), .C(_243_), .Y(_257_) );
OAI21X1 OAI21X1_41 ( .A(_184_), .B(_201_), .C(_257_), .Y(_258_) );
INVX1 INVX1_40 ( .A(_258_), .Y(_259_) );
NAND2X1 NAND2X1_32 ( .A(_129_), .B(_259_), .Y(_260_) );
INVX1 INVX1_41 ( .A(_184_), .Y(_261_) );
OAI21X1 OAI21X1_42 ( .A(_604_), .B(_227_), .C(_261_), .Y(_262_) );
AOI21X1 AOI21X1_21 ( .A(_262_), .B(_257_), .C(_129_), .Y(_263_) );
OAI21X1 OAI21X1_43 ( .A(_205_), .B(_240_), .C(_191_), .Y(_264_) );
NAND2X1 NAND2X1_33 ( .A(_198_), .B(_264_), .Y(_265_) );
NAND3X1 NAND3X1_44 ( .A(_527_), .B(_265_), .C(_243_), .Y(_266_) );
INVX1 INVX1_42 ( .A(_182_), .Y(_267_) );
OAI21X1 OAI21X1_44 ( .A(alu_inst_data_a_in_4_), .B(_267_), .C(_188_), .Y(_268_) );
OAI21X1 OAI21X1_45 ( .A(_604_), .B(_227_), .C(_268_), .Y(_269_) );
NAND3X1 NAND3X1_45 ( .A(_549_), .B(_266_), .C(_269_), .Y(_270_) );
OAI21X1 OAI21X1_46 ( .A(_270_), .B(_263_), .C(_260_), .Y(_271_) );
AOI21X1 AOI21X1_22 ( .A(_255_), .B(_271_), .C(_236_), .Y(_272_) );
INVX1 INVX1_43 ( .A(alu_inst_data_a_in_3_), .Y(_273_) );
NOR2X1 NOR2X1_17 ( .A(alu_inst_data_b_in_0_), .B(_273_), .Y(_274_) );
NOR2X1 NOR2X1_18 ( .A(_191_), .B(_274_), .Y(_275_) );
NAND3X1 NAND3X1_46 ( .A(_527_), .B(_275_), .C(_243_), .Y(_276_) );
OAI21X1 OAI21X1_47 ( .A(_604_), .B(_227_), .C(_273_), .Y(_277_) );
NAND3X1 NAND3X1_47 ( .A(_679_), .B(_276_), .C(_277_), .Y(_278_) );
AOI21X1 AOI21X1_23 ( .A(_277_), .B(_276_), .C(_679_), .Y(_279_) );
NOR2X1 NOR2X1_19 ( .A(alu_inst_data_a_in_2_), .B(_571_), .Y(_280_) );
OAI21X1 OAI21X1_48 ( .A(_280_), .B(_279_), .C(_278_), .Y(_281_) );
INVX1 INVX1_44 ( .A(_265_), .Y(_282_) );
NAND3X1 NAND3X1_48 ( .A(_527_), .B(_282_), .C(_243_), .Y(_283_) );
INVX1 INVX1_45 ( .A(_268_), .Y(_284_) );
OAI21X1 OAI21X1_49 ( .A(_604_), .B(_227_), .C(_284_), .Y(_285_) );
NAND3X1 NAND3X1_49 ( .A(alu_inst_data_b_in_2_), .B(_283_), .C(_285_), .Y(_286_) );
NAND2X1 NAND2X1_34 ( .A(_270_), .B(_286_), .Y(_287_) );
NAND3X1 NAND3X1_50 ( .A(alu_inst_data_b_in_3_), .B(_257_), .C(_262_), .Y(_288_) );
OAI21X1 OAI21X1_50 ( .A(_604_), .B(_227_), .C(_184_), .Y(_289_) );
XNOR2X1 XNOR2X1_5 ( .A(_206_), .B(_219_), .Y(_290_) );
NAND3X1 NAND3X1_51 ( .A(_527_), .B(_290_), .C(_243_), .Y(_291_) );
NAND3X1 NAND3X1_52 ( .A(_129_), .B(_291_), .C(_289_), .Y(_292_) );
AOI21X1 AOI21X1_24 ( .A(_288_), .B(_292_), .C(_287_), .Y(_293_) );
NAND3X1 NAND3X1_53 ( .A(_281_), .B(_293_), .C(_255_), .Y(_294_) );
AOI21X1 AOI21X1_25 ( .A(_272_), .B(_294_), .C(_225_), .Y(_295_) );
OAI21X1 OAI21X1_51 ( .A(_224_), .B(_295_), .C(_959_), .Y(_296_) );
INVX1 INVX1_46 ( .A(_296_), .Y(_297_) );
NAND2X1 NAND2X1_35 ( .A(alu_inst_data_b_in_6_), .B(_297_), .Y(_298_) );
NOR2X1 NOR2X1_20 ( .A(alu_inst_data_b_in_3_), .B(_258_), .Y(_299_) );
INVX1 INVX1_47 ( .A(_270_), .Y(_300_) );
NAND2X1 NAND2X1_36 ( .A(_288_), .B(_292_), .Y(_301_) );
AOI21X1 AOI21X1_26 ( .A(_300_), .B(_301_), .C(_299_), .Y(_302_) );
AND2X2 AND2X2_8 ( .A(_270_), .B(_286_), .Y(_303_) );
NAND3X1 NAND3X1_54 ( .A(_301_), .B(_303_), .C(_281_), .Y(_304_) );
AOI21X1 AOI21X1_27 ( .A(_304_), .B(_302_), .C(_254_), .Y(_305_) );
NAND3X1 NAND3X1_55 ( .A(_254_), .B(_302_), .C(_304_), .Y(_306_) );
INVX1 INVX1_48 ( .A(_306_), .Y(_307_) );
OAI21X1 OAI21X1_52 ( .A(_305_), .B(_307_), .C(_295_), .Y(_308_) );
OAI21X1 OAI21X1_53 ( .A(_251_), .B(_201_), .C(_231_), .Y(_309_) );
INVX1 INVX1_49 ( .A(_278_), .Y(_310_) );
OAI21X1 OAI21X1_54 ( .A(alu_inst_data_a_in_3_), .B(_201_), .C(_276_), .Y(_311_) );
NAND2X1 NAND2X1_37 ( .A(alu_inst_data_b_in_1_), .B(_311_), .Y(_312_) );
INVX1 INVX1_50 ( .A(_280_), .Y(_313_) );
AOI21X1 AOI21X1_28 ( .A(_312_), .B(_313_), .C(_310_), .Y(_314_) );
NAND3X1 NAND3X1_56 ( .A(_270_), .B(_286_), .C(_301_), .Y(_315_) );
OAI21X1 OAI21X1_55 ( .A(_315_), .B(_314_), .C(_302_), .Y(_316_) );
AOI21X1 AOI21X1_29 ( .A(_316_), .B(_255_), .C(_236_), .Y(_317_) );
OAI21X1 OAI21X1_56 ( .A(_225_), .B(_317_), .C(_309_), .Y(_318_) );
NAND3X1 NAND3X1_57 ( .A(_505_), .B(_318_), .C(_308_), .Y(_319_) );
OAI21X1 OAI21X1_57 ( .A(alu_inst_data_b_in_6_), .B(_297_), .C(_319_), .Y(_320_) );
XOR2X1 XOR2X1_3 ( .A(_296_), .B(_593_), .Y(_321_) );
INVX1 INVX1_51 ( .A(_305_), .Y(_322_) );
NAND3X1 NAND3X1_58 ( .A(_322_), .B(_306_), .C(_295_), .Y(_323_) );
OAI21X1 OAI21X1_58 ( .A(_238_), .B(_247_), .C(alu_inst_data_b_in_5_), .Y(_324_) );
AND2X2 AND2X2_9 ( .A(_253_), .B(_234_), .Y(_325_) );
NAND3X1 NAND3X1_59 ( .A(_229_), .B(_324_), .C(_325_), .Y(_326_) );
AOI21X1 AOI21X1_30 ( .A(_302_), .B(_304_), .C(_326_), .Y(_327_) );
OAI21X1 OAI21X1_59 ( .A(_236_), .B(_327_), .C(_516_), .Y(_328_) );
NAND3X1 NAND3X1_60 ( .A(_231_), .B(_233_), .C(_328_), .Y(_329_) );
NAND3X1 NAND3X1_61 ( .A(alu_inst_data_b_in_5_), .B(_323_), .C(_329_), .Y(_330_) );
AND2X2 AND2X2_10 ( .A(_330_), .B(_319_), .Y(_331_) );
AND2X2 AND2X2_11 ( .A(_331_), .B(_321_), .Y(_332_) );
AOI21X1 AOI21X1_31 ( .A(_281_), .B(_303_), .C(_300_), .Y(_333_) );
XOR2X1 XOR2X1_4 ( .A(_333_), .B(_301_), .Y(_334_) );
NAND2X1 NAND2X1_38 ( .A(_334_), .B(_295_), .Y(_335_) );
OAI21X1 OAI21X1_60 ( .A(_225_), .B(_317_), .C(_258_), .Y(_336_) );
NAND3X1 NAND3X1_62 ( .A(_152_), .B(_336_), .C(_335_), .Y(_337_) );
AOI21X1 AOI21X1_32 ( .A(_335_), .B(_336_), .C(_152_), .Y(_338_) );
NOR2X1 NOR2X1_21 ( .A(_287_), .B(_314_), .Y(_339_) );
NOR2X1 NOR2X1_22 ( .A(_303_), .B(_281_), .Y(_340_) );
OAI21X1 OAI21X1_61 ( .A(_339_), .B(_340_), .C(_295_), .Y(_341_) );
OAI21X1 OAI21X1_62 ( .A(_284_), .B(_201_), .C(_266_), .Y(_342_) );
OAI21X1 OAI21X1_63 ( .A(_225_), .B(_317_), .C(_342_), .Y(_343_) );
NAND3X1 NAND3X1_63 ( .A(_129_), .B(_343_), .C(_341_), .Y(_344_) );
OAI21X1 OAI21X1_64 ( .A(_344_), .B(_338_), .C(_337_), .Y(_345_) );
AOI22X1 AOI22X1_2 ( .A(_298_), .B(_320_), .C(_332_), .D(_345_), .Y(_346_) );
NOR2X1 NOR2X1_23 ( .A(alu_inst_data_a_in_1_), .B(_571_), .Y(_347_) );
INVX1 INVX1_52 ( .A(_236_), .Y(_348_) );
NAND2X1 NAND2X1_39 ( .A(_271_), .B(_255_), .Y(_349_) );
NAND3X1 NAND3X1_64 ( .A(_348_), .B(_349_), .C(_294_), .Y(_350_) );
NAND3X1 NAND3X1_65 ( .A(_278_), .B(_313_), .C(_312_), .Y(_351_) );
OAI21X1 OAI21X1_65 ( .A(_279_), .B(_310_), .C(_280_), .Y(_352_) );
NAND2X1 NAND2X1_40 ( .A(_351_), .B(_352_), .Y(_353_) );
INVX1 INVX1_53 ( .A(_353_), .Y(_354_) );
NAND3X1 NAND3X1_66 ( .A(_516_), .B(_354_), .C(_350_), .Y(_355_) );
INVX1 INVX1_54 ( .A(_311_), .Y(_356_) );
OAI21X1 OAI21X1_66 ( .A(_225_), .B(_317_), .C(_356_), .Y(_357_) );
AOI21X1 AOI21X1_33 ( .A(_357_), .B(_355_), .C(alu_inst_data_b_in_2_), .Y(_358_) );
NAND3X1 NAND3X1_67 ( .A(alu_inst_data_b_in_2_), .B(_355_), .C(_357_), .Y(_359_) );
INVX1 INVX1_55 ( .A(alu_inst_data_a_in_2_), .Y(_360_) );
NOR2X1 NOR2X1_24 ( .A(alu_inst_data_b_in_0_), .B(_360_), .Y(_361_) );
NOR2X1 NOR2X1_25 ( .A(_280_), .B(_361_), .Y(_362_) );
NAND3X1 NAND3X1_68 ( .A(_516_), .B(_362_), .C(_350_), .Y(_363_) );
OAI21X1 OAI21X1_67 ( .A(_225_), .B(_317_), .C(_360_), .Y(_364_) );
NAND3X1 NAND3X1_69 ( .A(_679_), .B(_363_), .C(_364_), .Y(_365_) );
INVX1 INVX1_56 ( .A(_365_), .Y(_366_) );
AOI21X1 AOI21X1_34 ( .A(_366_), .B(_359_), .C(_358_), .Y(_367_) );
OAI21X1 OAI21X1_68 ( .A(alu_inst_data_a_in_2_), .B(_295_), .C(_363_), .Y(_368_) );
NAND2X1 NAND2X1_41 ( .A(alu_inst_data_b_in_1_), .B(_368_), .Y(_369_) );
NAND3X1 NAND3X1_70 ( .A(_516_), .B(_353_), .C(_350_), .Y(_370_) );
OAI21X1 OAI21X1_69 ( .A(_225_), .B(_317_), .C(_311_), .Y(_371_) );
NAND3X1 NAND3X1_71 ( .A(alu_inst_data_b_in_2_), .B(_370_), .C(_371_), .Y(_372_) );
NAND3X1 NAND3X1_72 ( .A(_549_), .B(_355_), .C(_357_), .Y(_373_) );
NAND2X1 NAND2X1_42 ( .A(_372_), .B(_373_), .Y(_374_) );
NAND3X1 NAND3X1_73 ( .A(_365_), .B(_369_), .C(_374_), .Y(_375_) );
OAI21X1 OAI21X1_70 ( .A(_347_), .B(_375_), .C(_367_), .Y(_376_) );
NAND3X1 NAND3X1_74 ( .A(alu_inst_data_b_in_4_), .B(_336_), .C(_335_), .Y(_377_) );
OAI21X1 OAI21X1_71 ( .A(_259_), .B(_295_), .C(_335_), .Y(_378_) );
NAND2X1 NAND2X1_43 ( .A(_152_), .B(_378_), .Y(_379_) );
NOR2X1 NOR2X1_26 ( .A(_340_), .B(_339_), .Y(_380_) );
NAND2X1 NAND2X1_44 ( .A(_380_), .B(_295_), .Y(_381_) );
INVX1 INVX1_57 ( .A(_342_), .Y(_382_) );
OAI21X1 OAI21X1_72 ( .A(_225_), .B(_317_), .C(_382_), .Y(_383_) );
NAND3X1 NAND3X1_75 ( .A(alu_inst_data_b_in_3_), .B(_383_), .C(_381_), .Y(_384_) );
NAND2X1 NAND2X1_45 ( .A(_384_), .B(_344_), .Y(_385_) );
AOI21X1 AOI21X1_35 ( .A(_377_), .B(_379_), .C(_385_), .Y(_386_) );
NAND3X1 NAND3X1_76 ( .A(_332_), .B(_386_), .C(_376_), .Y(_387_) );
NAND2X1 NAND2X1_46 ( .A(_346_), .B(_387_), .Y(_388_) );
INVX1 INVX1_58 ( .A(_321_), .Y(_389_) );
INVX1 INVX1_59 ( .A(_345_), .Y(_390_) );
AOI21X1 AOI21X1_36 ( .A(_364_), .B(_363_), .C(_679_), .Y(_391_) );
OAI21X1 OAI21X1_73 ( .A(_347_), .B(_391_), .C(_365_), .Y(_392_) );
AOI21X1 AOI21X1_37 ( .A(_392_), .B(_359_), .C(_358_), .Y(_393_) );
INVX1 INVX1_60 ( .A(_338_), .Y(_394_) );
AND2X2 AND2X2_12 ( .A(_344_), .B(_384_), .Y(_395_) );
NAND3X1 NAND3X1_77 ( .A(_337_), .B(_394_), .C(_395_), .Y(_396_) );
OAI21X1 OAI21X1_74 ( .A(_396_), .B(_393_), .C(_390_), .Y(_397_) );
NAND2X1 NAND2X1_47 ( .A(_331_), .B(_397_), .Y(_398_) );
AOI21X1 AOI21X1_38 ( .A(_398_), .B(_319_), .C(_389_), .Y(_399_) );
INVX1 INVX1_61 ( .A(_319_), .Y(_400_) );
INVX1 INVX1_62 ( .A(_331_), .Y(_401_) );
INVX1 INVX1_63 ( .A(_358_), .Y(_402_) );
INVX1 INVX1_64 ( .A(_347_), .Y(_403_) );
NAND3X1 NAND3X1_78 ( .A(_365_), .B(_403_), .C(_369_), .Y(_404_) );
NAND3X1 NAND3X1_79 ( .A(_402_), .B(_365_), .C(_404_), .Y(_405_) );
NAND3X1 NAND3X1_80 ( .A(_359_), .B(_386_), .C(_405_), .Y(_407_) );
AOI21X1 AOI21X1_39 ( .A(_407_), .B(_390_), .C(_401_), .Y(_408_) );
NOR3X1 NOR3X1_2 ( .A(_400_), .B(_321_), .C(_408_), .Y(_409_) );
OAI21X1 OAI21X1_75 ( .A(_399_), .B(_409_), .C(_388_), .Y(_410_) );
OAI21X1 OAI21X1_76 ( .A(_593_), .B(_296_), .C(_320_), .Y(_411_) );
NAND2X1 NAND2X1_48 ( .A(_321_), .B(_331_), .Y(_412_) );
OAI21X1 OAI21X1_77 ( .A(_390_), .B(_412_), .C(_411_), .Y(_413_) );
NOR2X1 NOR2X1_27 ( .A(_396_), .B(_412_), .Y(_414_) );
AOI21X1 AOI21X1_40 ( .A(_414_), .B(_376_), .C(_413_), .Y(_415_) );
AOI21X1 AOI21X1_41 ( .A(_415_), .B(_297_), .C(alu_inst_data_b_in_7_), .Y(_416_) );
NAND2X1 NAND2X1_49 ( .A(_416_), .B(_410_), .Y(_418_) );
NOR2X1 NOR2X1_28 ( .A(alu_inst_data_a_in_7_), .B(_582_), .Y(_419_) );
AOI21X1 AOI21X1_42 ( .A(_387_), .B(_346_), .C(alu_inst_data_b_in_7_), .Y(_420_) );
NOR2X1 NOR2X1_29 ( .A(_331_), .B(_397_), .Y(_421_) );
OAI21X1 OAI21X1_78 ( .A(_408_), .B(_421_), .C(_420_), .Y(_422_) );
NAND2X1 NAND2X1_50 ( .A(_318_), .B(_308_), .Y(_423_) );
OAI21X1 OAI21X1_79 ( .A(alu_inst_data_b_in_7_), .B(_415_), .C(_423_), .Y(_424_) );
NAND3X1 NAND3X1_81 ( .A(_593_), .B(_424_), .C(_422_), .Y(_425_) );
OR2X2 OR2X2_1 ( .A(_425_), .B(_419_), .Y(_426_) );
AOI22X1 AOI22X1_3 ( .A(alu_inst_data_b_in_7_), .B(_560_), .C(_410_), .D(_416_), .Y(_427_) );
NAND3X1 NAND3X1_82 ( .A(_401_), .B(_390_), .C(_407_), .Y(_429_) );
NAND3X1 NAND3X1_83 ( .A(_398_), .B(_429_), .C(_420_), .Y(_430_) );
INVX1 INVX1_65 ( .A(_423_), .Y(_431_) );
OAI21X1 OAI21X1_80 ( .A(alu_inst_data_b_in_7_), .B(_415_), .C(_431_), .Y(_432_) );
NAND3X1 NAND3X1_84 ( .A(alu_inst_data_b_in_6_), .B(_432_), .C(_430_), .Y(_433_) );
AND2X2 AND2X2_13 ( .A(_425_), .B(_433_), .Y(_434_) );
NAND2X1 NAND2X1_51 ( .A(_377_), .B(_379_), .Y(_435_) );
OAI21X1 OAI21X1_81 ( .A(_385_), .B(_393_), .C(_344_), .Y(_436_) );
NOR2X1 NOR2X1_30 ( .A(_435_), .B(_436_), .Y(_437_) );
AND2X2 AND2X2_14 ( .A(_436_), .B(_435_), .Y(_438_) );
OAI21X1 OAI21X1_82 ( .A(_437_), .B(_438_), .C(_420_), .Y(_440_) );
OAI21X1 OAI21X1_83 ( .A(alu_inst_data_b_in_7_), .B(_415_), .C(_378_), .Y(_441_) );
AOI21X1 AOI21X1_43 ( .A(_440_), .B(_441_), .C(_505_), .Y(_442_) );
NAND3X1 NAND3X1_85 ( .A(_505_), .B(_441_), .C(_440_), .Y(_443_) );
XOR2X1 XOR2X1_5 ( .A(_393_), .B(_395_), .Y(_444_) );
NAND3X1 NAND3X1_86 ( .A(_582_), .B(_444_), .C(_388_), .Y(_445_) );
OAI21X1 OAI21X1_84 ( .A(_328_), .B(_380_), .C(_343_), .Y(_446_) );
OAI21X1 OAI21X1_85 ( .A(alu_inst_data_b_in_7_), .B(_415_), .C(_446_), .Y(_447_) );
NAND3X1 NAND3X1_87 ( .A(_152_), .B(_445_), .C(_447_), .Y(_448_) );
AOI21X1 AOI21X1_44 ( .A(_443_), .B(_448_), .C(_442_), .Y(_449_) );
NAND3X1 NAND3X1_88 ( .A(_434_), .B(_427_), .C(_449_), .Y(_451_) );
NAND3X1 NAND3X1_89 ( .A(_418_), .B(_426_), .C(_451_), .Y(_452_) );
NOR2X1 NOR2X1_31 ( .A(alu_inst_data_a_in_0_), .B(_571_), .Y(_453_) );
OAI21X1 OAI21X1_86 ( .A(_311_), .B(_295_), .C(_355_), .Y(_454_) );
INVX1 INVX1_66 ( .A(_454_), .Y(_455_) );
XOR2X1 XOR2X1_6 ( .A(_392_), .B(_374_), .Y(_456_) );
NAND2X1 NAND2X1_52 ( .A(_456_), .B(_420_), .Y(_457_) );
OAI21X1 OAI21X1_87 ( .A(_455_), .B(_420_), .C(_457_), .Y(_458_) );
AOI22X1 AOI22X1_4 ( .A(alu_inst_data_b_in_1_), .B(_453_), .C(_458_), .D(_129_), .Y(_459_) );
INVX1 INVX1_67 ( .A(_404_), .Y(_460_) );
AOI21X1 AOI21X1_45 ( .A(_369_), .B(_365_), .C(_403_), .Y(_462_) );
OAI21X1 OAI21X1_88 ( .A(_460_), .B(_462_), .C(_420_), .Y(_463_) );
OAI21X1 OAI21X1_89 ( .A(alu_inst_data_b_in_7_), .B(_415_), .C(_368_), .Y(_464_) );
NAND3X1 NAND3X1_90 ( .A(_549_), .B(_464_), .C(_463_), .Y(_465_) );
INVX1 INVX1_68 ( .A(_368_), .Y(_466_) );
OAI21X1 OAI21X1_90 ( .A(alu_inst_data_b_in_7_), .B(_415_), .C(_466_), .Y(_467_) );
NOR2X1 NOR2X1_32 ( .A(_462_), .B(_460_), .Y(_468_) );
NAND2X1 NAND2X1_53 ( .A(_468_), .B(_420_), .Y(_469_) );
NAND3X1 NAND3X1_91 ( .A(alu_inst_data_b_in_2_), .B(_467_), .C(_469_), .Y(_470_) );
AND2X2 AND2X2_15 ( .A(_465_), .B(_470_), .Y(_471_) );
MUX2X1 MUX2X1_1 ( .A(_456_), .B(_454_), .S(_420_), .Y(_473_) );
NAND2X1 NAND2X1_54 ( .A(_582_), .B(_388_), .Y(_474_) );
OAI21X1 OAI21X1_91 ( .A(_571_), .B(_474_), .C(alu_inst_data_a_in_1_), .Y(_475_) );
INVX1 INVX1_69 ( .A(_453_), .Y(_476_) );
AOI22X1 AOI22X1_5 ( .A(_679_), .B(_476_), .C(_420_), .D(_347_), .Y(_477_) );
AOI22X1 AOI22X1_6 ( .A(_475_), .B(_477_), .C(_473_), .D(alu_inst_data_b_in_3_), .Y(_478_) );
NAND3X1 NAND3X1_92 ( .A(_459_), .B(_478_), .C(_471_), .Y(_479_) );
OAI21X1 OAI21X1_92 ( .A(alu_inst_data_b_in_3_), .B(_473_), .C(_465_), .Y(_480_) );
OAI21X1 OAI21X1_93 ( .A(_129_), .B(_458_), .C(_480_), .Y(_481_) );
NAND3X1 NAND3X1_93 ( .A(alu_inst_data_b_in_5_), .B(_441_), .C(_440_), .Y(_482_) );
INVX1 INVX1_70 ( .A(_378_), .Y(_484_) );
OAI21X1 OAI21X1_94 ( .A(alu_inst_data_b_in_7_), .B(_415_), .C(_484_), .Y(_485_) );
INVX1 INVX1_71 ( .A(_435_), .Y(_486_) );
NOR2X1 NOR2X1_33 ( .A(_486_), .B(_436_), .Y(_487_) );
AND2X2 AND2X2_16 ( .A(_436_), .B(_486_), .Y(_488_) );
OAI21X1 OAI21X1_95 ( .A(_487_), .B(_488_), .C(_420_), .Y(_489_) );
NAND3X1 NAND3X1_94 ( .A(_505_), .B(_485_), .C(_489_), .Y(_490_) );
NAND3X1 NAND3X1_95 ( .A(alu_inst_data_b_in_4_), .B(_445_), .C(_447_), .Y(_491_) );
XOR2X1 XOR2X1_7 ( .A(_393_), .B(_385_), .Y(_492_) );
NAND3X1 NAND3X1_96 ( .A(_582_), .B(_492_), .C(_388_), .Y(_493_) );
INVX1 INVX1_72 ( .A(_446_), .Y(_495_) );
OAI21X1 OAI21X1_96 ( .A(alu_inst_data_b_in_7_), .B(_415_), .C(_495_), .Y(_496_) );
NAND3X1 NAND3X1_97 ( .A(_152_), .B(_493_), .C(_496_), .Y(_497_) );
AOI22X1 AOI22X1_7 ( .A(_491_), .B(_497_), .C(_490_), .D(_482_), .Y(_498_) );
NAND3X1 NAND3X1_98 ( .A(_498_), .B(_434_), .C(_427_), .Y(_499_) );
AOI21X1 AOI21X1_46 ( .A(_479_), .B(_481_), .C(_499_), .Y(_500_) );
OAI21X1 OAI21X1_97 ( .A(_452_), .B(_500_), .C(_483_), .Y(_501_) );
NOR2X1 NOR2X1_34 ( .A(alu_inst_data_b_in_7_), .B(_560_), .Y(_502_) );
INVX1 INVX1_73 ( .A(_502_), .Y(_503_) );
INVX1 INVX1_74 ( .A(alu_inst_data_a_in_6_), .Y(_504_) );
NOR2X1 NOR2X1_35 ( .A(_593_), .B(_504_), .Y(_506_) );
NOR2X1 NOR2X1_36 ( .A(alu_inst_data_b_in_6_), .B(alu_inst_data_a_in_6_), .Y(_507_) );
NOR2X1 NOR2X1_37 ( .A(_505_), .B(_818_), .Y(_508_) );
NOR2X1 NOR2X1_38 ( .A(alu_inst_data_b_in_5_), .B(alu_inst_data_a_in_5_), .Y(_509_) );
INVX1 INVX1_75 ( .A(alu_inst_data_a_in_1_), .Y(_510_) );
NOR2X1 NOR2X1_39 ( .A(_510_), .B(_679_), .Y(_511_) );
NOR2X1 NOR2X1_40 ( .A(alu_inst_data_a_in_1_), .B(alu_inst_data_b_in_1_), .Y(_512_) );
OAI21X1 OAI21X1_98 ( .A(_511_), .B(_512_), .C(_476_), .Y(_513_) );
OAI21X1 OAI21X1_99 ( .A(_510_), .B(alu_inst_data_b_in_1_), .C(_513_), .Y(_514_) );
NOR2X1 NOR2X1_41 ( .A(_549_), .B(_360_), .Y(_515_) );
NOR2X1 NOR2X1_42 ( .A(alu_inst_data_b_in_2_), .B(alu_inst_data_a_in_2_), .Y(_517_) );
OAI21X1 OAI21X1_100 ( .A(_515_), .B(_517_), .C(_514_), .Y(_518_) );
OAI21X1 OAI21X1_101 ( .A(alu_inst_data_b_in_2_), .B(_360_), .C(_518_), .Y(_519_) );
OAI21X1 OAI21X1_102 ( .A(_129_), .B(alu_inst_data_a_in_3_), .C(_519_), .Y(_520_) );
OAI21X1 OAI21X1_103 ( .A(alu_inst_data_b_in_3_), .B(_273_), .C(_520_), .Y(_521_) );
NOR2X1 NOR2X1_43 ( .A(_152_), .B(_840_), .Y(_522_) );
NOR2X1 NOR2X1_44 ( .A(alu_inst_data_b_in_4_), .B(alu_inst_data_a_in_4_), .Y(_523_) );
OAI21X1 OAI21X1_104 ( .A(_522_), .B(_523_), .C(_521_), .Y(_524_) );
OAI21X1 OAI21X1_105 ( .A(alu_inst_data_b_in_4_), .B(_840_), .C(_524_), .Y(_525_) );
OAI21X1 OAI21X1_106 ( .A(_508_), .B(_509_), .C(_525_), .Y(_526_) );
OAI21X1 OAI21X1_107 ( .A(alu_inst_data_b_in_5_), .B(_818_), .C(_526_), .Y(_528_) );
OAI21X1 OAI21X1_108 ( .A(_506_), .B(_507_), .C(_528_), .Y(_529_) );
OAI21X1 OAI21X1_109 ( .A(alu_inst_data_b_in_6_), .B(_504_), .C(_529_), .Y(_530_) );
INVX1 INVX1_76 ( .A(_530_), .Y(_531_) );
OAI21X1 OAI21X1_110 ( .A(_419_), .B(_531_), .C(_503_), .Y(_532_) );
INVX1 INVX1_77 ( .A(alu_inst_alu_func_in_2_), .Y(_533_) );
INVX1 INVX1_78 ( .A(alu_inst_alu_func_in_3_), .Y(_534_) );
NOR2X1 NOR2X1_45 ( .A(_533_), .B(_534_), .Y(_535_) );
NOR2X1 NOR2X1_46 ( .A(alu_inst_alu_func_in_1_), .B(alu_inst_alu_func_in_0_), .Y(_536_) );
NAND2X1 NAND2X1_55 ( .A(_536_), .B(_535_), .Y(_537_) );
NOR2X1 NOR2X1_47 ( .A(_537_), .B(_532_), .Y(_539_) );
NOR2X1 NOR2X1_48 ( .A(_509_), .B(_508_), .Y(_540_) );
INVX1 INVX1_79 ( .A(_540_), .Y(_541_) );
OAI21X1 OAI21X1_111 ( .A(_522_), .B(_523_), .C(_541_), .Y(_542_) );
NOR2X1 NOR2X1_49 ( .A(_582_), .B(_560_), .Y(_543_) );
NOR2X1 NOR2X1_50 ( .A(_507_), .B(_506_), .Y(_544_) );
INVX1 INVX1_80 ( .A(_544_), .Y(_545_) );
NOR2X1 NOR2X1_51 ( .A(alu_inst_data_b_in_7_), .B(alu_inst_data_a_in_7_), .Y(_546_) );
OAI21X1 OAI21X1_112 ( .A(_543_), .B(_546_), .C(_545_), .Y(_547_) );
NOR2X1 NOR2X1_52 ( .A(_542_), .B(_547_), .Y(_548_) );
INVX1 INVX1_81 ( .A(_548_), .Y(_550_) );
NOR2X1 NOR2X1_53 ( .A(_517_), .B(_515_), .Y(_551_) );
INVX1 INVX1_82 ( .A(_551_), .Y(_552_) );
NOR2X1 NOR2X1_54 ( .A(_129_), .B(_273_), .Y(_553_) );
NOR2X1 NOR2X1_55 ( .A(alu_inst_data_b_in_3_), .B(alu_inst_data_a_in_3_), .Y(_554_) );
OAI21X1 OAI21X1_113 ( .A(_553_), .B(_554_), .C(_552_), .Y(_555_) );
NOR2X1 NOR2X1_56 ( .A(_512_), .B(_511_), .Y(_556_) );
INVX1 INVX1_83 ( .A(_556_), .Y(_557_) );
INVX1 INVX1_84 ( .A(alu_inst_data_a_in_0_), .Y(_558_) );
NOR2X1 NOR2X1_57 ( .A(_571_), .B(_558_), .Y(_559_) );
NOR2X1 NOR2X1_58 ( .A(alu_inst_data_b_in_0_), .B(alu_inst_data_a_in_0_), .Y(_561_) );
OAI21X1 OAI21X1_114 ( .A(_559_), .B(_561_), .C(_557_), .Y(_562_) );
OR2X2 OR2X2_2 ( .A(_555_), .B(_562_), .Y(_563_) );
NOR2X1 NOR2X1_59 ( .A(_563_), .B(_550_), .Y(_564_) );
INVX1 INVX1_85 ( .A(_564_), .Y(_565_) );
NOR2X1 NOR2X1_60 ( .A(alu_inst_alu_func_in_2_), .B(_534_), .Y(_566_) );
NOR2X1 NOR2X1_61 ( .A(alu_inst_alu_func_in_0_), .B(_417_), .Y(_567_) );
NAND2X1 NAND2X1_56 ( .A(_566_), .B(_567_), .Y(_568_) );
NOR2X1 NOR2X1_62 ( .A(alu_inst_alu_func_in_1_), .B(_428_), .Y(_569_) );
INVX1 INVX1_86 ( .A(_569_), .Y(_570_) );
NOR2X1 NOR2X1_63 ( .A(alu_inst_alu_func_in_3_), .B(_533_), .Y(_572_) );
INVX1 INVX1_87 ( .A(_572_), .Y(_573_) );
NOR2X1 NOR2X1_64 ( .A(_570_), .B(_573_), .Y(_574_) );
INVX1 INVX1_88 ( .A(_574_), .Y(_575_) );
NOR2X1 NOR2X1_65 ( .A(_561_), .B(_559_), .Y(_576_) );
INVX1 INVX1_89 ( .A(_536_), .Y(_577_) );
INVX1 INVX1_90 ( .A(_566_), .Y(_578_) );
NOR2X1 NOR2X1_66 ( .A(_577_), .B(_578_), .Y(_579_) );
NOR2X1 NOR2X1_67 ( .A(alu_inst_alu_func_in_1_), .B(_472_), .Y(_580_) );
OAI21X1 OAI21X1_115 ( .A(_580_), .B(_579_), .C(_576_), .Y(_581_) );
OAI21X1 OAI21X1_116 ( .A(_561_), .B(_575_), .C(_581_), .Y(_583_) );
INVX1 INVX1_91 ( .A(_559_), .Y(_584_) );
INVX1 INVX1_92 ( .A(_567_), .Y(_585_) );
OAI21X1 OAI21X1_117 ( .A(_585_), .B(_573_), .C(_584_), .Y(_586_) );
NOR2X1 NOR2X1_68 ( .A(_577_), .B(_573_), .Y(_587_) );
OAI21X1 OAI21X1_118 ( .A(_584_), .B(_587_), .C(_586_), .Y(_588_) );
NOR2X1 NOR2X1_69 ( .A(_578_), .B(_570_), .Y(_589_) );
INVX1 INVX1_93 ( .A(_589_), .Y(_590_) );
NOR2X1 NOR2X1_70 ( .A(_472_), .B(_585_), .Y(_591_) );
INVX1 INVX1_94 ( .A(_591_), .Y(_592_) );
OAI21X1 OAI21X1_119 ( .A(_584_), .B(_592_), .C(_590_), .Y(_594_) );
OAI21X1 OAI21X1_120 ( .A(_559_), .B(_561_), .C(_594_), .Y(_595_) );
INVX1 INVX1_95 ( .A(_535_), .Y(_596_) );
NOR2X1 NOR2X1_71 ( .A(_570_), .B(_596_), .Y(_597_) );
NOR2X1 NOR2X1_72 ( .A(_573_), .B(_450_), .Y(_598_) );
AOI22X1 AOI22X1_8 ( .A(_597_), .B(alu_inst_data_a_in_1_), .C(_561_), .D(_598_), .Y(_599_) );
NAND3X1 NAND3X1_99 ( .A(_588_), .B(_595_), .C(_599_), .Y(_600_) );
NOR2X1 NOR2X1_73 ( .A(_583_), .B(_600_), .Y(_601_) );
OAI21X1 OAI21X1_121 ( .A(_568_), .B(_565_), .C(_601_), .Y(_602_) );
NOR2X1 NOR2X1_74 ( .A(_602_), .B(_539_), .Y(_603_) );
AOI21X1 AOI21X1_47 ( .A(_501_), .B(_603_), .C(_406_), .Y(alu_inst_alu_out_comp_0_) );
INVX1 INVX1_96 ( .A(_483_), .Y(_605_) );
NOR2X1 NOR2X1_75 ( .A(_578_), .B(_450_), .Y(_606_) );
AND2X2 AND2X2_17 ( .A(_532_), .B(_565_), .Y(_607_) );
NOR2X1 NOR2X1_76 ( .A(_472_), .B(_570_), .Y(_608_) );
INVX1 INVX1_97 ( .A(_608_), .Y(_609_) );
NAND2X1 NAND2X1_57 ( .A(_453_), .B(_556_), .Y(_610_) );
NAND2X1 NAND2X1_58 ( .A(_513_), .B(_610_), .Y(_611_) );
INVX1 INVX1_98 ( .A(_511_), .Y(_612_) );
INVX1 INVX1_99 ( .A(_587_), .Y(_613_) );
OAI21X1 OAI21X1_122 ( .A(_612_), .B(_613_), .C(_590_), .Y(_615_) );
OAI21X1 OAI21X1_123 ( .A(_511_), .B(_512_), .C(_615_), .Y(_616_) );
OAI21X1 OAI21X1_124 ( .A(_512_), .B(_575_), .C(_616_), .Y(_617_) );
NAND2X1 NAND2X1_59 ( .A(_461_), .B(_536_), .Y(_618_) );
NOR2X1 NOR2X1_77 ( .A(_584_), .B(_557_), .Y(_619_) );
NOR2X1 NOR2X1_78 ( .A(_618_), .B(_619_), .Y(_620_) );
OAI21X1 OAI21X1_125 ( .A(_556_), .B(_559_), .C(_620_), .Y(_621_) );
NOR2X1 NOR2X1_79 ( .A(_585_), .B(_573_), .Y(_622_) );
OAI21X1 OAI21X1_126 ( .A(_510_), .B(_679_), .C(_622_), .Y(_623_) );
INVX1 INVX1_100 ( .A(_579_), .Y(_624_) );
NOR2X1 NOR2X1_80 ( .A(_585_), .B(_596_), .Y(_626_) );
INVX1 INVX1_101 ( .A(_626_), .Y(_627_) );
OAI22X1 OAI22X1_1 ( .A(_557_), .B(_624_), .C(_558_), .D(_627_), .Y(_628_) );
NAND2X1 NAND2X1_60 ( .A(alu_inst_data_a_in_1_), .B(alu_inst_data_b_in_0_), .Y(_629_) );
OAI21X1 OAI21X1_127 ( .A(_679_), .B(_558_), .C(_629_), .Y(_630_) );
OAI21X1 OAI21X1_128 ( .A(_612_), .B(_584_), .C(_630_), .Y(_631_) );
AOI22X1 AOI22X1_9 ( .A(_597_), .B(alu_inst_data_a_in_2_), .C(_512_), .D(_598_), .Y(_632_) );
OAI21X1 OAI21X1_129 ( .A(_592_), .B(_631_), .C(_632_), .Y(_633_) );
NOR2X1 NOR2X1_81 ( .A(_628_), .B(_633_), .Y(_634_) );
NAND3X1 NAND3X1_100 ( .A(_623_), .B(_621_), .C(_634_), .Y(_635_) );
NOR2X1 NOR2X1_82 ( .A(_617_), .B(_635_), .Y(_637_) );
OAI21X1 OAI21X1_130 ( .A(_609_), .B(_611_), .C(_637_), .Y(_638_) );
OR2X2 OR2X2_3 ( .A(_539_), .B(_638_), .Y(_639_) );
AOI21X1 AOI21X1_48 ( .A(_606_), .B(_607_), .C(_639_), .Y(_640_) );
OAI21X1 OAI21X1_131 ( .A(_605_), .B(_474_), .C(_640_), .Y(_641_) );
AND2X2 AND2X2_18 ( .A(_641_), .B(alu_inst_alu_out_comp_valid), .Y(alu_inst_alu_out_comp_1_) );
NOR2X1 NOR2X1_83 ( .A(_612_), .B(_584_), .Y(_642_) );
NAND2X1 NAND2X1_61 ( .A(alu_inst_data_a_in_2_), .B(alu_inst_data_b_in_1_), .Y(_643_) );
NAND2X1 NAND2X1_62 ( .A(alu_inst_data_a_in_2_), .B(alu_inst_data_b_in_0_), .Y(_644_) );
OAI21X1 OAI21X1_132 ( .A(_510_), .B(_679_), .C(_644_), .Y(_645_) );
OAI21X1 OAI21X1_133 ( .A(_629_), .B(_643_), .C(_645_), .Y(_647_) );
OAI21X1 OAI21X1_134 ( .A(_549_), .B(_558_), .C(_647_), .Y(_648_) );
INVX1 INVX1_102 ( .A(_647_), .Y(_649_) );
NAND3X1 NAND3X1_101 ( .A(alu_inst_data_b_in_2_), .B(alu_inst_data_a_in_0_), .C(_649_), .Y(_650_) );
AND2X2 AND2X2_19 ( .A(_650_), .B(_648_), .Y(_651_) );
NAND2X1 NAND2X1_63 ( .A(_642_), .B(_651_), .Y(_652_) );
INVX1 INVX1_103 ( .A(_652_), .Y(_653_) );
OAI21X1 OAI21X1_135 ( .A(_642_), .B(_651_), .C(_591_), .Y(_654_) );
NOR2X1 NOR2X1_84 ( .A(_654_), .B(_653_), .Y(_655_) );
OAI21X1 OAI21X1_136 ( .A(_511_), .B(_619_), .C(_551_), .Y(_656_) );
INVX1 INVX1_104 ( .A(_656_), .Y(_658_) );
NOR2X1 NOR2X1_85 ( .A(_472_), .B(_577_), .Y(_659_) );
OAI21X1 OAI21X1_137 ( .A(_512_), .B(_584_), .C(_612_), .Y(_660_) );
OAI21X1 OAI21X1_138 ( .A(_551_), .B(_660_), .C(_659_), .Y(_661_) );
NOR2X1 NOR2X1_86 ( .A(_661_), .B(_658_), .Y(_662_) );
AOI21X1 AOI21X1_49 ( .A(_514_), .B(_552_), .C(_609_), .Y(_663_) );
OAI21X1 OAI21X1_139 ( .A(_514_), .B(_552_), .C(_663_), .Y(_664_) );
OAI21X1 OAI21X1_140 ( .A(_515_), .B(_624_), .C(_575_), .Y(_665_) );
OAI21X1 OAI21X1_141 ( .A(alu_inst_data_b_in_2_), .B(alu_inst_data_a_in_2_), .C(_665_), .Y(_666_) );
INVX1 INVX1_105 ( .A(_622_), .Y(_667_) );
AOI22X1 AOI22X1_10 ( .A(_597_), .B(alu_inst_data_a_in_3_), .C(alu_inst_data_a_in_1_), .D(_626_), .Y(_669_) );
OAI21X1 OAI21X1_142 ( .A(_515_), .B(_667_), .C(_669_), .Y(_670_) );
INVX1 INVX1_106 ( .A(_515_), .Y(_671_) );
OAI21X1 OAI21X1_143 ( .A(_578_), .B(_570_), .C(_613_), .Y(_672_) );
INVX1 INVX1_107 ( .A(_672_), .Y(_673_) );
OAI21X1 OAI21X1_144 ( .A(_589_), .B(_598_), .C(_517_), .Y(_674_) );
OAI21X1 OAI21X1_145 ( .A(_671_), .B(_673_), .C(_674_), .Y(_675_) );
NOR2X1 NOR2X1_87 ( .A(_670_), .B(_675_), .Y(_676_) );
NAND3X1 NAND3X1_102 ( .A(_664_), .B(_666_), .C(_676_), .Y(_677_) );
OR2X2 OR2X2_4 ( .A(_677_), .B(_662_), .Y(_678_) );
NOR2X1 NOR2X1_88 ( .A(_655_), .B(_678_), .Y(_680_) );
OAI21X1 OAI21X1_146 ( .A(_605_), .B(_328_), .C(_680_), .Y(_681_) );
AND2X2 AND2X2_20 ( .A(_681_), .B(alu_inst_alu_out_comp_valid), .Y(alu_inst_alu_out_comp_2_) );
NOR2X1 NOR2X1_89 ( .A(_129_), .B(_558_), .Y(_682_) );
OAI21X1 OAI21X1_147 ( .A(_612_), .B(_644_), .C(_650_), .Y(_683_) );
NAND2X1 NAND2X1_64 ( .A(alu_inst_data_a_in_3_), .B(alu_inst_data_b_in_1_), .Y(_684_) );
OAI21X1 OAI21X1_148 ( .A(_273_), .B(_571_), .C(_643_), .Y(_685_) );
OAI21X1 OAI21X1_149 ( .A(_644_), .B(_684_), .C(_685_), .Y(_686_) );
OAI21X1 OAI21X1_150 ( .A(_510_), .B(_549_), .C(_686_), .Y(_687_) );
NAND2X1 NAND2X1_65 ( .A(alu_inst_data_a_in_1_), .B(alu_inst_data_b_in_2_), .Y(_688_) );
OR2X2 OR2X2_5 ( .A(_686_), .B(_688_), .Y(_690_) );
AND2X2 AND2X2_21 ( .A(_690_), .B(_687_), .Y(_691_) );
NOR2X1 NOR2X1_90 ( .A(_683_), .B(_691_), .Y(_692_) );
NAND2X1 NAND2X1_66 ( .A(_683_), .B(_691_), .Y(_693_) );
INVX1 INVX1_108 ( .A(_693_), .Y(_694_) );
NOR2X1 NOR2X1_91 ( .A(_692_), .B(_694_), .Y(_695_) );
XOR2X1 XOR2X1_8 ( .A(_695_), .B(_682_), .Y(_696_) );
OR2X2 OR2X2_6 ( .A(_696_), .B(_653_), .Y(_697_) );
NAND2X1 NAND2X1_67 ( .A(_653_), .B(_696_), .Y(_698_) );
INVX1 INVX1_109 ( .A(_698_), .Y(_699_) );
NOR2X1 NOR2X1_92 ( .A(_592_), .B(_699_), .Y(_701_) );
INVX1 INVX1_110 ( .A(_554_), .Y(_702_) );
OAI21X1 OAI21X1_151 ( .A(_549_), .B(_360_), .C(_656_), .Y(_703_) );
INVX1 INVX1_111 ( .A(_703_), .Y(_704_) );
AOI22X1 AOI22X1_11 ( .A(_519_), .B(_608_), .C(_704_), .D(_659_), .Y(_705_) );
NOR2X1 NOR2X1_93 ( .A(_553_), .B(_705_), .Y(_706_) );
OAI21X1 OAI21X1_152 ( .A(_553_), .B(_624_), .C(_575_), .Y(_707_) );
OAI21X1 OAI21X1_153 ( .A(_707_), .B(_706_), .C(_702_), .Y(_708_) );
OAI22X1 OAI22X1_2 ( .A(_519_), .B(_609_), .C(_618_), .D(_704_), .Y(_709_) );
OAI21X1 OAI21X1_154 ( .A(_553_), .B(_554_), .C(_709_), .Y(_710_) );
INVX1 INVX1_112 ( .A(_553_), .Y(_712_) );
AOI22X1 AOI22X1_12 ( .A(_622_), .B(_712_), .C(alu_inst_data_a_in_4_), .D(_597_), .Y(_713_) );
OAI21X1 OAI21X1_155 ( .A(_360_), .B(_627_), .C(_713_), .Y(_714_) );
OAI21X1 OAI21X1_156 ( .A(_589_), .B(_598_), .C(_554_), .Y(_715_) );
OAI21X1 OAI21X1_157 ( .A(_712_), .B(_673_), .C(_715_), .Y(_716_) );
NOR2X1 NOR2X1_94 ( .A(_714_), .B(_716_), .Y(_717_) );
NAND3X1 NAND3X1_103 ( .A(_710_), .B(_717_), .C(_708_), .Y(_718_) );
AOI21X1 AOI21X1_50 ( .A(_701_), .B(_697_), .C(_718_), .Y(_719_) );
OAI21X1 OAI21X1_158 ( .A(_605_), .B(_244_), .C(_719_), .Y(_720_) );
AND2X2 AND2X2_22 ( .A(_720_), .B(alu_inst_alu_out_comp_valid), .Y(alu_inst_alu_out_comp_3_) );
INVX1 INVX1_113 ( .A(_682_), .Y(_722_) );
OAI21X1 OAI21X1_159 ( .A(_722_), .B(_692_), .C(_693_), .Y(_723_) );
NOR2X1 NOR2X1_95 ( .A(_510_), .B(_152_), .Y(_724_) );
INVX1 INVX1_114 ( .A(_724_), .Y(_725_) );
OAI22X1 OAI22X1_3 ( .A(_510_), .B(_129_), .C(_152_), .D(_558_), .Y(_726_) );
OAI21X1 OAI21X1_160 ( .A(_722_), .B(_725_), .C(_726_), .Y(_727_) );
OAI21X1 OAI21X1_161 ( .A(_644_), .B(_684_), .C(_690_), .Y(_728_) );
XOR2X1 XOR2X1_9 ( .A(_851_), .B(_684_), .Y(_729_) );
OR2X2 OR2X2_7 ( .A(_729_), .B(_671_), .Y(_730_) );
OAI21X1 OAI21X1_162 ( .A(_549_), .B(_360_), .C(_729_), .Y(_731_) );
AND2X2 AND2X2_23 ( .A(_730_), .B(_731_), .Y(_733_) );
NOR2X1 NOR2X1_96 ( .A(_728_), .B(_733_), .Y(_734_) );
NAND2X1 NAND2X1_68 ( .A(_728_), .B(_733_), .Y(_735_) );
INVX1 INVX1_115 ( .A(_735_), .Y(_736_) );
NOR2X1 NOR2X1_97 ( .A(_734_), .B(_736_), .Y(_737_) );
XNOR2X1 XNOR2X1_6 ( .A(_737_), .B(_727_), .Y(_738_) );
NAND2X1 NAND2X1_69 ( .A(_723_), .B(_738_), .Y(_739_) );
INVX1 INVX1_116 ( .A(_739_), .Y(_740_) );
NOR2X1 NOR2X1_98 ( .A(_723_), .B(_738_), .Y(_741_) );
NOR2X1 NOR2X1_99 ( .A(_741_), .B(_740_), .Y(_742_) );
AOI21X1 AOI21X1_51 ( .A(_742_), .B(_699_), .C(_592_), .Y(_744_) );
OAI21X1 OAI21X1_163 ( .A(_699_), .B(_742_), .C(_744_), .Y(_745_) );
NOR2X1 NOR2X1_100 ( .A(_523_), .B(_522_), .Y(_746_) );
INVX1 INVX1_117 ( .A(_746_), .Y(_747_) );
AOI21X1 AOI21X1_52 ( .A(_521_), .B(_747_), .C(_609_), .Y(_748_) );
OAI21X1 OAI21X1_164 ( .A(_521_), .B(_747_), .C(_748_), .Y(_749_) );
OAI21X1 OAI21X1_165 ( .A(_554_), .B(_704_), .C(_712_), .Y(_750_) );
INVX1 INVX1_118 ( .A(_750_), .Y(_751_) );
AOI21X1 AOI21X1_53 ( .A(_751_), .B(_747_), .C(_618_), .Y(_752_) );
OAI21X1 OAI21X1_166 ( .A(_747_), .B(_751_), .C(_752_), .Y(_753_) );
INVX1 INVX1_119 ( .A(_522_), .Y(_755_) );
OAI21X1 OAI21X1_167 ( .A(_523_), .B(_624_), .C(_667_), .Y(_756_) );
AOI22X1 AOI22X1_13 ( .A(_597_), .B(alu_inst_data_a_in_5_), .C(alu_inst_data_a_in_3_), .D(_626_), .Y(_757_) );
OAI21X1 OAI21X1_168 ( .A(alu_inst_data_b_in_4_), .B(alu_inst_data_a_in_4_), .C(_574_), .Y(_758_) );
OAI21X1 OAI21X1_169 ( .A(_450_), .B(_573_), .C(_590_), .Y(_759_) );
AOI22X1 AOI22X1_14 ( .A(_672_), .B(_522_), .C(_523_), .D(_759_), .Y(_760_) );
NAND3X1 NAND3X1_104 ( .A(_757_), .B(_758_), .C(_760_), .Y(_761_) );
AOI21X1 AOI21X1_54 ( .A(_755_), .B(_756_), .C(_761_), .Y(_762_) );
NAND3X1 NAND3X1_105 ( .A(_749_), .B(_762_), .C(_753_), .Y(_763_) );
AOI21X1 AOI21X1_55 ( .A(_267_), .B(_483_), .C(_763_), .Y(_764_) );
AOI21X1 AOI21X1_56 ( .A(_764_), .B(_745_), .C(_406_), .Y(alu_inst_alu_out_comp_4_) );
NAND2X1 NAND2X1_70 ( .A(_699_), .B(_742_), .Y(_766_) );
NOR2X1 NOR2X1_101 ( .A(_722_), .B(_725_), .Y(_767_) );
OAI21X1 OAI21X1_170 ( .A(_727_), .B(_734_), .C(_735_), .Y(_768_) );
NOR2X1 NOR2X1_102 ( .A(_505_), .B(_558_), .Y(_769_) );
NAND2X1 NAND2X1_71 ( .A(alu_inst_data_b_in_3_), .B(alu_inst_data_a_in_2_), .Y(_770_) );
XNOR2X1 XNOR2X1_7 ( .A(_724_), .B(_770_), .Y(_771_) );
XOR2X1 XOR2X1_10 ( .A(_771_), .B(_769_), .Y(_772_) );
OAI21X1 OAI21X1_171 ( .A(_862_), .B(_684_), .C(_730_), .Y(_773_) );
NAND2X1 NAND2X1_72 ( .A(alu_inst_data_a_in_5_), .B(alu_inst_data_b_in_1_), .Y(_774_) );
NAND2X1 NAND2X1_73 ( .A(alu_inst_data_a_in_4_), .B(alu_inst_data_b_in_1_), .Y(_776_) );
OAI21X1 OAI21X1_172 ( .A(_818_), .B(_571_), .C(_776_), .Y(_777_) );
OAI21X1 OAI21X1_173 ( .A(_774_), .B(_862_), .C(_777_), .Y(_778_) );
OAI21X1 OAI21X1_174 ( .A(_273_), .B(_549_), .C(_778_), .Y(_779_) );
NAND2X1 NAND2X1_74 ( .A(alu_inst_data_a_in_3_), .B(alu_inst_data_b_in_2_), .Y(_780_) );
OR2X2 OR2X2_8 ( .A(_778_), .B(_780_), .Y(_781_) );
AND2X2 AND2X2_24 ( .A(_781_), .B(_779_), .Y(_782_) );
XOR2X1 XOR2X1_11 ( .A(_782_), .B(_773_), .Y(_783_) );
XOR2X1 XOR2X1_12 ( .A(_783_), .B(_772_), .Y(_784_) );
XOR2X1 XOR2X1_13 ( .A(_784_), .B(_768_), .Y(_785_) );
OR2X2 OR2X2_9 ( .A(_785_), .B(_767_), .Y(_787_) );
NAND2X1 NAND2X1_75 ( .A(_767_), .B(_785_), .Y(_788_) );
NAND2X1 NAND2X1_76 ( .A(_788_), .B(_787_), .Y(_789_) );
INVX1 INVX1_120 ( .A(_789_), .Y(_790_) );
NOR2X1 NOR2X1_103 ( .A(_740_), .B(_790_), .Y(_791_) );
NAND2X1 NAND2X1_77 ( .A(_740_), .B(_790_), .Y(_792_) );
INVX1 INVX1_121 ( .A(_792_), .Y(_793_) );
OAI21X1 OAI21X1_175 ( .A(_791_), .B(_793_), .C(_766_), .Y(_794_) );
NOR2X1 NOR2X1_104 ( .A(_789_), .B(_766_), .Y(_795_) );
NOR2X1 NOR2X1_105 ( .A(_592_), .B(_795_), .Y(_796_) );
AOI21X1 AOI21X1_57 ( .A(_525_), .B(_541_), .C(_609_), .Y(_798_) );
OAI21X1 OAI21X1_176 ( .A(_541_), .B(_525_), .C(_798_), .Y(_799_) );
OAI21X1 OAI21X1_177 ( .A(_523_), .B(_751_), .C(_755_), .Y(_800_) );
NOR2X1 NOR2X1_106 ( .A(_747_), .B(_751_), .Y(_801_) );
OAI21X1 OAI21X1_178 ( .A(_522_), .B(_801_), .C(_540_), .Y(_802_) );
INVX1 INVX1_122 ( .A(_802_), .Y(_803_) );
NOR2X1 NOR2X1_107 ( .A(_618_), .B(_803_), .Y(_804_) );
OAI21X1 OAI21X1_179 ( .A(_540_), .B(_800_), .C(_804_), .Y(_805_) );
OAI21X1 OAI21X1_180 ( .A(_505_), .B(_818_), .C(_579_), .Y(_806_) );
AOI21X1 AOI21X1_58 ( .A(_806_), .B(_575_), .C(_509_), .Y(_807_) );
AOI22X1 AOI22X1_15 ( .A(_597_), .B(alu_inst_data_a_in_6_), .C(alu_inst_data_a_in_4_), .D(_626_), .Y(_809_) );
OAI21X1 OAI21X1_181 ( .A(_505_), .B(_818_), .C(_622_), .Y(_810_) );
AOI22X1 AOI22X1_16 ( .A(_672_), .B(_508_), .C(_509_), .D(_759_), .Y(_811_) );
NAND3X1 NAND3X1_106 ( .A(_809_), .B(_810_), .C(_811_), .Y(_812_) );
NOR2X1 NOR2X1_108 ( .A(_807_), .B(_812_), .Y(_813_) );
NAND3X1 NAND3X1_107 ( .A(_799_), .B(_813_), .C(_805_), .Y(_814_) );
AOI21X1 AOI21X1_59 ( .A(_794_), .B(_796_), .C(_814_), .Y(_815_) );
OAI21X1 OAI21X1_182 ( .A(_605_), .B(_1003_), .C(_815_), .Y(_816_) );
AND2X2 AND2X2_25 ( .A(_816_), .B(alu_inst_alu_out_comp_valid), .Y(alu_inst_alu_out_comp_5_) );
AOI21X1 AOI21X1_60 ( .A(_528_), .B(_545_), .C(_609_), .Y(_817_) );
OAI21X1 OAI21X1_183 ( .A(_545_), .B(_528_), .C(_817_), .Y(_819_) );
NAND2X1 NAND2X1_78 ( .A(_768_), .B(_784_), .Y(_820_) );
NAND2X1 NAND2X1_79 ( .A(_820_), .B(_788_), .Y(_821_) );
NOR2X1 NOR2X1_109 ( .A(_593_), .B(_558_), .Y(_822_) );
NAND2X1 NAND2X1_80 ( .A(_769_), .B(_771_), .Y(_823_) );
OAI21X1 OAI21X1_184 ( .A(_725_), .B(_770_), .C(_823_), .Y(_824_) );
NOR2X1 NOR2X1_110 ( .A(_822_), .B(_824_), .Y(_825_) );
NAND2X1 NAND2X1_81 ( .A(_822_), .B(_824_), .Y(_826_) );
INVX1 INVX1_123 ( .A(_826_), .Y(_827_) );
NOR2X1 NOR2X1_111 ( .A(_825_), .B(_827_), .Y(_828_) );
NAND2X1 NAND2X1_82 ( .A(_773_), .B(_782_), .Y(_830_) );
NAND2X1 NAND2X1_83 ( .A(_772_), .B(_783_), .Y(_831_) );
NAND2X1 NAND2X1_84 ( .A(_830_), .B(_831_), .Y(_832_) );
NOR2X1 NOR2X1_112 ( .A(_510_), .B(_505_), .Y(_833_) );
NAND2X1 NAND2X1_85 ( .A(alu_inst_data_b_in_4_), .B(alu_inst_data_a_in_2_), .Y(_834_) );
XNOR2X1 XNOR2X1_8 ( .A(_553_), .B(_834_), .Y(_835_) );
XOR2X1 XOR2X1_14 ( .A(_835_), .B(_833_), .Y(_836_) );
NOR2X1 NOR2X1_113 ( .A(_818_), .B(_571_), .Y(_837_) );
INVX1 INVX1_124 ( .A(_837_), .Y(_838_) );
OAI21X1 OAI21X1_185 ( .A(_838_), .B(_776_), .C(_781_), .Y(_839_) );
NOR2X1 NOR2X1_114 ( .A(_504_), .B(_679_), .Y(_841_) );
INVX1 INVX1_125 ( .A(_841_), .Y(_842_) );
OAI21X1 OAI21X1_186 ( .A(_504_), .B(_571_), .C(_774_), .Y(_843_) );
OAI21X1 OAI21X1_187 ( .A(_838_), .B(_842_), .C(_843_), .Y(_844_) );
OAI21X1 OAI21X1_188 ( .A(_840_), .B(_549_), .C(_844_), .Y(_845_) );
NAND2X1 NAND2X1_86 ( .A(alu_inst_data_a_in_4_), .B(alu_inst_data_b_in_2_), .Y(_846_) );
OR2X2 OR2X2_10 ( .A(_844_), .B(_846_), .Y(_847_) );
AND2X2 AND2X2_26 ( .A(_847_), .B(_845_), .Y(_848_) );
XOR2X1 XOR2X1_15 ( .A(_848_), .B(_839_), .Y(_849_) );
XOR2X1 XOR2X1_16 ( .A(_849_), .B(_836_), .Y(_850_) );
NOR2X1 NOR2X1_115 ( .A(_832_), .B(_850_), .Y(_852_) );
NAND2X1 NAND2X1_87 ( .A(_832_), .B(_850_), .Y(_853_) );
INVX1 INVX1_126 ( .A(_853_), .Y(_854_) );
NOR2X1 NOR2X1_116 ( .A(_852_), .B(_854_), .Y(_855_) );
XOR2X1 XOR2X1_17 ( .A(_855_), .B(_828_), .Y(_856_) );
NAND2X1 NAND2X1_88 ( .A(_821_), .B(_856_), .Y(_857_) );
INVX1 INVX1_127 ( .A(_857_), .Y(_858_) );
NOR2X1 NOR2X1_117 ( .A(_821_), .B(_856_), .Y(_859_) );
NOR2X1 NOR2X1_118 ( .A(_859_), .B(_858_), .Y(_860_) );
NOR2X1 NOR2X1_119 ( .A(_793_), .B(_860_), .Y(_861_) );
INVX1 INVX1_128 ( .A(_860_), .Y(_863_) );
NOR2X1 NOR2X1_120 ( .A(_792_), .B(_863_), .Y(_864_) );
NOR2X1 NOR2X1_121 ( .A(_861_), .B(_864_), .Y(_865_) );
NAND2X1 NAND2X1_89 ( .A(_795_), .B(_865_), .Y(_866_) );
INVX1 INVX1_129 ( .A(_866_), .Y(_867_) );
OAI21X1 OAI21X1_189 ( .A(_795_), .B(_865_), .C(_591_), .Y(_868_) );
NOR2X1 NOR2X1_122 ( .A(_868_), .B(_867_), .Y(_869_) );
NOR2X1 NOR2X1_123 ( .A(_508_), .B(_803_), .Y(_870_) );
AOI21X1 AOI21X1_61 ( .A(_870_), .B(_545_), .C(_618_), .Y(_871_) );
OAI21X1 OAI21X1_190 ( .A(_545_), .B(_870_), .C(_871_), .Y(_872_) );
AND2X2 AND2X2_27 ( .A(_765_), .B(_775_), .Y(_874_) );
OAI21X1 OAI21X1_191 ( .A(_507_), .B(_624_), .C(_667_), .Y(_875_) );
OAI21X1 OAI21X1_192 ( .A(_593_), .B(_504_), .C(_875_), .Y(_876_) );
INVX1 INVX1_130 ( .A(_507_), .Y(_877_) );
NAND2X1 NAND2X1_90 ( .A(alu_inst_data_a_in_7_), .B(_597_), .Y(_878_) );
OAI21X1 OAI21X1_193 ( .A(_818_), .B(_627_), .C(_878_), .Y(_879_) );
AOI21X1 AOI21X1_62 ( .A(_877_), .B(_574_), .C(_879_), .Y(_880_) );
AOI22X1 AOI22X1_17 ( .A(_672_), .B(_506_), .C(_507_), .D(_759_), .Y(_881_) );
NAND3X1 NAND3X1_108 ( .A(_876_), .B(_881_), .C(_880_), .Y(_882_) );
AOI21X1 AOI21X1_63 ( .A(_874_), .B(_483_), .C(_882_), .Y(_883_) );
NAND2X1 NAND2X1_91 ( .A(_883_), .B(_872_), .Y(_885_) );
NOR2X1 NOR2X1_124 ( .A(_885_), .B(_869_), .Y(_886_) );
AOI21X1 AOI21X1_64 ( .A(_886_), .B(_819_), .C(_406_), .Y(alu_inst_alu_out_comp_6_) );
OAI21X1 OAI21X1_194 ( .A(_792_), .B(_863_), .C(_866_), .Y(_887_) );
INVX1 INVX1_131 ( .A(_828_), .Y(_888_) );
OAI21X1 OAI21X1_195 ( .A(_888_), .B(_852_), .C(_853_), .Y(_889_) );
NOR2X1 NOR2X1_125 ( .A(_510_), .B(_593_), .Y(_890_) );
NAND2X1 NAND2X1_92 ( .A(_833_), .B(_835_), .Y(_891_) );
OAI21X1 OAI21X1_196 ( .A(_712_), .B(_834_), .C(_891_), .Y(_892_) );
XOR2X1 XOR2X1_18 ( .A(_892_), .B(_890_), .Y(_893_) );
INVX1 INVX1_132 ( .A(_893_), .Y(_895_) );
OAI21X1 OAI21X1_197 ( .A(_582_), .B(_558_), .C(_895_), .Y(_896_) );
NAND3X1 NAND3X1_109 ( .A(alu_inst_data_b_in_7_), .B(alu_inst_data_a_in_0_), .C(_893_), .Y(_897_) );
AND2X2 AND2X2_28 ( .A(_896_), .B(_897_), .Y(_898_) );
NAND2X1 NAND2X1_93 ( .A(_839_), .B(_848_), .Y(_899_) );
NAND2X1 NAND2X1_94 ( .A(_836_), .B(_849_), .Y(_900_) );
NAND2X1 NAND2X1_95 ( .A(_899_), .B(_900_), .Y(_901_) );
NOR2X1 NOR2X1_126 ( .A(_505_), .B(_360_), .Y(_902_) );
AOI22X1 AOI22X1_18 ( .A(alu_inst_data_b_in_4_), .B(alu_inst_data_a_in_3_), .C(alu_inst_data_a_in_4_), .D(alu_inst_data_b_in_3_), .Y(_903_) );
AOI21X1 AOI21X1_65 ( .A(_553_), .B(_522_), .C(_903_), .Y(_904_) );
XOR2X1 XOR2X1_19 ( .A(_904_), .B(_902_), .Y(_906_) );
OAI21X1 OAI21X1_198 ( .A(_838_), .B(_842_), .C(_847_), .Y(_907_) );
NOR2X1 NOR2X1_127 ( .A(_818_), .B(_549_), .Y(_908_) );
INVX1 INVX1_133 ( .A(_908_), .Y(_909_) );
NOR2X1 NOR2X1_128 ( .A(_560_), .B(_571_), .Y(_910_) );
INVX1 INVX1_134 ( .A(_910_), .Y(_911_) );
NOR2X1 NOR2X1_129 ( .A(_911_), .B(_842_), .Y(_912_) );
OAI21X1 OAI21X1_199 ( .A(_560_), .B(_571_), .C(_842_), .Y(_913_) );
INVX1 INVX1_135 ( .A(_913_), .Y(_914_) );
OAI21X1 OAI21X1_200 ( .A(_912_), .B(_914_), .C(_909_), .Y(_915_) );
INVX1 INVX1_136 ( .A(_912_), .Y(_917_) );
NAND3X1 NAND3X1_110 ( .A(_908_), .B(_913_), .C(_917_), .Y(_918_) );
AND2X2 AND2X2_29 ( .A(_918_), .B(_915_), .Y(_919_) );
XOR2X1 XOR2X1_20 ( .A(_919_), .B(_907_), .Y(_920_) );
XOR2X1 XOR2X1_21 ( .A(_920_), .B(_906_), .Y(_921_) );
XOR2X1 XOR2X1_22 ( .A(_921_), .B(_901_), .Y(_922_) );
XOR2X1 XOR2X1_23 ( .A(_922_), .B(_898_), .Y(_923_) );
NOR2X1 NOR2X1_130 ( .A(_889_), .B(_923_), .Y(_924_) );
NAND2X1 NAND2X1_96 ( .A(_889_), .B(_923_), .Y(_925_) );
INVX1 INVX1_137 ( .A(_925_), .Y(_926_) );
NOR2X1 NOR2X1_131 ( .A(_924_), .B(_926_), .Y(_928_) );
XOR2X1 XOR2X1_24 ( .A(_928_), .B(_827_), .Y(_929_) );
XOR2X1 XOR2X1_25 ( .A(_929_), .B(_858_), .Y(_930_) );
AOI21X1 AOI21X1_66 ( .A(_887_), .B(_930_), .C(_592_), .Y(_931_) );
OAI21X1 OAI21X1_201 ( .A(_887_), .B(_930_), .C(_931_), .Y(_932_) );
NOR2X1 NOR2X1_132 ( .A(_546_), .B(_543_), .Y(_933_) );
OAI21X1 OAI21X1_202 ( .A(_933_), .B(_531_), .C(_608_), .Y(_934_) );
AOI21X1 AOI21X1_67 ( .A(_531_), .B(_933_), .C(_934_), .Y(_935_) );
INVX1 INVX1_138 ( .A(_933_), .Y(_936_) );
OAI21X1 OAI21X1_203 ( .A(_508_), .B(_803_), .C(_544_), .Y(_937_) );
OAI21X1 OAI21X1_204 ( .A(_593_), .B(_504_), .C(_937_), .Y(_939_) );
INVX1 INVX1_139 ( .A(_939_), .Y(_940_) );
NOR2X1 NOR2X1_133 ( .A(_936_), .B(_940_), .Y(_941_) );
OAI21X1 OAI21X1_205 ( .A(_933_), .B(_939_), .C(_659_), .Y(_942_) );
OAI21X1 OAI21X1_206 ( .A(_543_), .B(_546_), .C(_589_), .Y(_943_) );
OAI21X1 OAI21X1_207 ( .A(_936_), .B(_624_), .C(_943_), .Y(_944_) );
INVX1 INVX1_140 ( .A(_625_), .Y(_945_) );
NAND2X1 NAND2X1_97 ( .A(_527_), .B(_945_), .Y(_946_) );
OAI21X1 OAI21X1_208 ( .A(alu_inst_data_a_in_7_), .B(_571_), .C(_483_), .Y(_947_) );
OAI22X1 OAI22X1_4 ( .A(_543_), .B(_667_), .C(_546_), .D(_575_), .Y(_948_) );
NAND2X1 NAND2X1_98 ( .A(_546_), .B(_598_), .Y(_950_) );
OAI21X1 OAI21X1_209 ( .A(_504_), .B(_627_), .C(_950_), .Y(_951_) );
NOR2X1 NOR2X1_134 ( .A(_951_), .B(_948_), .Y(_952_) );
OAI21X1 OAI21X1_210 ( .A(_946_), .B(_947_), .C(_952_), .Y(_953_) );
OR2X2 OR2X2_11 ( .A(_953_), .B(_944_), .Y(_954_) );
AOI21X1 AOI21X1_68 ( .A(_543_), .B(_587_), .C(_954_), .Y(_955_) );
OAI21X1 OAI21X1_211 ( .A(_942_), .B(_941_), .C(_955_), .Y(_956_) );
NOR2X1 NOR2X1_135 ( .A(_935_), .B(_956_), .Y(_957_) );
AOI21X1 AOI21X1_69 ( .A(_932_), .B(_957_), .C(_406_), .Y(alu_inst_alu_out_comp_7_) );
INVX1 INVX1_141 ( .A(_929_), .Y(_958_) );
OAI21X1 OAI21X1_212 ( .A(_864_), .B(_867_), .C(_930_), .Y(_960_) );
OAI21X1 OAI21X1_213 ( .A(_857_), .B(_958_), .C(_960_), .Y(_961_) );
OAI21X1 OAI21X1_214 ( .A(_826_), .B(_924_), .C(_925_), .Y(_962_) );
NAND2X1 NAND2X1_99 ( .A(_890_), .B(_892_), .Y(_963_) );
NAND2X1 NAND2X1_100 ( .A(_963_), .B(_897_), .Y(_964_) );
NAND2X1 NAND2X1_101 ( .A(_901_), .B(_921_), .Y(_965_) );
NAND2X1 NAND2X1_102 ( .A(_898_), .B(_922_), .Y(_966_) );
NAND2X1 NAND2X1_103 ( .A(_965_), .B(_966_), .Y(_967_) );
NOR2X1 NOR2X1_136 ( .A(_593_), .B(_360_), .Y(_968_) );
NAND2X1 NAND2X1_104 ( .A(_902_), .B(_904_), .Y(_969_) );
OAI21X1 OAI21X1_215 ( .A(_712_), .B(_755_), .C(_969_), .Y(_971_) );
XOR2X1 XOR2X1_26 ( .A(_971_), .B(_968_), .Y(_972_) );
INVX1 INVX1_142 ( .A(_972_), .Y(_973_) );
OAI21X1 OAI21X1_216 ( .A(_510_), .B(_582_), .C(_973_), .Y(_974_) );
NAND3X1 NAND3X1_111 ( .A(alu_inst_data_a_in_1_), .B(alu_inst_data_b_in_7_), .C(_972_), .Y(_975_) );
AND2X2 AND2X2_30 ( .A(_974_), .B(_975_), .Y(_976_) );
NAND2X1 NAND2X1_105 ( .A(_907_), .B(_919_), .Y(_977_) );
NAND2X1 NAND2X1_106 ( .A(_906_), .B(_920_), .Y(_978_) );
NAND2X1 NAND2X1_107 ( .A(_977_), .B(_978_), .Y(_979_) );
NOR2X1 NOR2X1_137 ( .A(_505_), .B(_273_), .Y(_980_) );
NAND2X1 NAND2X1_108 ( .A(alu_inst_data_a_in_5_), .B(alu_inst_data_b_in_3_), .Y(_982_) );
XNOR2X1 XNOR2X1_9 ( .A(_522_), .B(_982_), .Y(_983_) );
XOR2X1 XOR2X1_27 ( .A(_983_), .B(_980_), .Y(_984_) );
OAI21X1 OAI21X1_217 ( .A(_909_), .B(_914_), .C(_917_), .Y(_985_) );
INVX1 INVX1_143 ( .A(_985_), .Y(_986_) );
INVX1 INVX1_144 ( .A(_646_), .Y(_987_) );
NOR2X1 NOR2X1_138 ( .A(_679_), .B(_987_), .Y(_988_) );
NAND3X1 NAND3X1_112 ( .A(alu_inst_data_a_in_6_), .B(alu_inst_data_b_in_2_), .C(_988_), .Y(_989_) );
INVX1 INVX1_145 ( .A(_988_), .Y(_990_) );
OAI21X1 OAI21X1_218 ( .A(_504_), .B(_549_), .C(_990_), .Y(_991_) );
NAND2X1 NAND2X1_109 ( .A(_989_), .B(_991_), .Y(_993_) );
XOR2X1 XOR2X1_28 ( .A(_993_), .B(_986_), .Y(_994_) );
XOR2X1 XOR2X1_29 ( .A(_994_), .B(_984_), .Y(_995_) );
NOR2X1 NOR2X1_139 ( .A(_979_), .B(_995_), .Y(_996_) );
NAND2X1 NAND2X1_110 ( .A(_979_), .B(_995_), .Y(_997_) );
INVX1 INVX1_146 ( .A(_997_), .Y(_998_) );
NOR2X1 NOR2X1_140 ( .A(_996_), .B(_998_), .Y(_999_) );
NOR2X1 NOR2X1_141 ( .A(_976_), .B(_999_), .Y(_1000_) );
NAND2X1 NAND2X1_111 ( .A(_976_), .B(_999_), .Y(_1001_) );
INVX1 INVX1_147 ( .A(_1001_), .Y(_1002_) );
NOR2X1 NOR2X1_142 ( .A(_1000_), .B(_1002_), .Y(_1004_) );
XNOR2X1 XNOR2X1_10 ( .A(_1004_), .B(_967_), .Y(_1005_) );
XNOR2X1 XNOR2X1_11 ( .A(_1005_), .B(_964_), .Y(_1006_) );
XOR2X1 XOR2X1_30 ( .A(_1006_), .B(_962_), .Y(_1007_) );
NAND2X1 NAND2X1_112 ( .A(_1007_), .B(_961_), .Y(_1008_) );
OR2X2 OR2X2_12 ( .A(_961_), .B(_1007_), .Y(_1009_) );
NAND3X1 NAND3X1_113 ( .A(_591_), .B(_1008_), .C(_1009_), .Y(_1010_) );
INVX1 INVX1_148 ( .A(_543_), .Y(_1011_) );
OAI21X1 OAI21X1_219 ( .A(_546_), .B(_940_), .C(_1011_), .Y(_1012_) );
AOI22X1 AOI22X1_19 ( .A(alu_inst_data_a_in_7_), .B(_626_), .C(_1012_), .D(_659_), .Y(_1013_) );
INVX1 INVX1_149 ( .A(_532_), .Y(_1015_) );
NAND2X1 NAND2X1_113 ( .A(_571_), .B(_483_), .Y(_1016_) );
AOI21X1 AOI21X1_70 ( .A(alu_inst_alu_func_in_1_), .B(_572_), .C(_589_), .Y(_1017_) );
OAI21X1 OAI21X1_220 ( .A(_946_), .B(_1016_), .C(_1017_), .Y(_1018_) );
AOI21X1 AOI21X1_71 ( .A(_1015_), .B(_608_), .C(_1018_), .Y(_1019_) );
AND2X2 AND2X2_31 ( .A(_1013_), .B(_1019_), .Y(_1020_) );
AOI21X1 AOI21X1_72 ( .A(_1010_), .B(_1020_), .C(_406_), .Y(alu_inst_alu_out_comp_8_) );
NAND2X1 NAND2X1_114 ( .A(_962_), .B(_1006_), .Y(_1021_) );
NAND2X1 NAND2X1_115 ( .A(_1021_), .B(_1008_), .Y(_1022_) );
NAND2X1 NAND2X1_116 ( .A(_967_), .B(_1004_), .Y(_1023_) );
INVX1 INVX1_150 ( .A(_1005_), .Y(_1025_) );
NAND2X1 NAND2X1_117 ( .A(_964_), .B(_1025_), .Y(_1026_) );
NAND2X1 NAND2X1_118 ( .A(_1023_), .B(_1026_), .Y(_1027_) );
NAND2X1 NAND2X1_119 ( .A(_968_), .B(_971_), .Y(_1028_) );
NAND2X1 NAND2X1_120 ( .A(_1028_), .B(_975_), .Y(_1029_) );
NOR2X1 NOR2X1_143 ( .A(_998_), .B(_1002_), .Y(_1030_) );
NOR2X1 NOR2X1_144 ( .A(_593_), .B(_273_), .Y(_1031_) );
NAND2X1 NAND2X1_121 ( .A(_980_), .B(_983_), .Y(_1032_) );
OAI21X1 OAI21X1_221 ( .A(_755_), .B(_982_), .C(_1032_), .Y(_1033_) );
XOR2X1 XOR2X1_31 ( .A(_1033_), .B(_1031_), .Y(_1034_) );
INVX1 INVX1_151 ( .A(_1034_), .Y(_1036_) );
OAI21X1 OAI21X1_222 ( .A(_582_), .B(_360_), .C(_1036_), .Y(_1037_) );
NAND3X1 NAND3X1_114 ( .A(alu_inst_data_b_in_7_), .B(alu_inst_data_a_in_2_), .C(_1034_), .Y(_1038_) );
AND2X2 AND2X2_32 ( .A(_1037_), .B(_1038_), .Y(_1039_) );
NAND2X1 NAND2X1_122 ( .A(_984_), .B(_994_), .Y(_1040_) );
OAI21X1 OAI21X1_223 ( .A(_986_), .B(_993_), .C(_1040_), .Y(_1041_) );
NOR2X1 NOR2X1_145 ( .A(_505_), .B(_840_), .Y(_1042_) );
NOR2X1 NOR2X1_146 ( .A(_504_), .B(_152_), .Y(_1043_) );
INVX1 INVX1_152 ( .A(_1043_), .Y(_1044_) );
NOR2X1 NOR2X1_147 ( .A(_982_), .B(_1044_), .Y(_1045_) );
AOI22X1 AOI22X1_20 ( .A(alu_inst_data_a_in_6_), .B(alu_inst_data_b_in_3_), .C(alu_inst_data_a_in_5_), .D(alu_inst_data_b_in_4_), .Y(_1047_) );
NOR2X1 NOR2X1_148 ( .A(_1047_), .B(_1045_), .Y(_1048_) );
XNOR2X1 XNOR2X1_12 ( .A(_1048_), .B(_1042_), .Y(_1049_) );
NAND3X1 NAND3X1_115 ( .A(alu_inst_data_b_in_2_), .B(_842_), .C(_646_), .Y(_1050_) );
XOR2X1 XOR2X1_32 ( .A(_1049_), .B(_1050_), .Y(_1051_) );
XOR2X1 XOR2X1_33 ( .A(_1041_), .B(_1051_), .Y(_1052_) );
XNOR2X1 XNOR2X1_13 ( .A(_1052_), .B(_1039_), .Y(_1053_) );
XOR2X1 XOR2X1_34 ( .A(_1030_), .B(_1053_), .Y(_1054_) );
XNOR2X1 XNOR2X1_14 ( .A(_1054_), .B(_1029_), .Y(_1055_) );
XNOR2X1 XNOR2X1_15 ( .A(_1027_), .B(_1055_), .Y(_1056_) );
NAND2X1 NAND2X1_123 ( .A(_1056_), .B(_1022_), .Y(_1058_) );
OR2X2 OR2X2_13 ( .A(_1022_), .B(_1056_), .Y(_1059_) );
NAND3X1 NAND3X1_116 ( .A(_591_), .B(_1058_), .C(_1059_), .Y(_1060_) );
AOI21X1 AOI21X1_73 ( .A(_1060_), .B(_1019_), .C(_406_), .Y(alu_inst_alu_out_comp_9_) );
INVX1 INVX1_153 ( .A(_1027_), .Y(_1061_) );
OAI21X1 OAI21X1_224 ( .A(_1061_), .B(_1055_), .C(_1058_), .Y(_1062_) );
NAND2X1 NAND2X1_124 ( .A(_1029_), .B(_1054_), .Y(_1063_) );
OAI21X1 OAI21X1_225 ( .A(_1030_), .B(_1053_), .C(_1063_), .Y(_1064_) );
NAND2X1 NAND2X1_125 ( .A(_1031_), .B(_1033_), .Y(_1065_) );
NAND2X1 NAND2X1_126 ( .A(_1065_), .B(_1038_), .Y(_1066_) );
INVX1 INVX1_154 ( .A(_1066_), .Y(_0_) );
NAND2X1 NAND2X1_127 ( .A(_1051_), .B(_1041_), .Y(_1_) );
NAND2X1 NAND2X1_128 ( .A(_1039_), .B(_1052_), .Y(_2_) );
NAND2X1 NAND2X1_129 ( .A(_1_), .B(_2_), .Y(_3_) );
NOR2X1 NOR2X1_149 ( .A(_582_), .B(_273_), .Y(_4_) );
NOR2X1 NOR2X1_150 ( .A(_593_), .B(_840_), .Y(_5_) );
NAND2X1 NAND2X1_130 ( .A(_1042_), .B(_1048_), .Y(_6_) );
OAI21X1 OAI21X1_226 ( .A(_982_), .B(_1044_), .C(_6_), .Y(_7_) );
XOR2X1 XOR2X1_35 ( .A(_7_), .B(_5_), .Y(_8_) );
XOR2X1 XOR2X1_36 ( .A(_8_), .B(_4_), .Y(_9_) );
OAI21X1 OAI21X1_227 ( .A(_1050_), .B(_1049_), .C(_989_), .Y(_11_) );
XOR2X1 XOR2X1_37 ( .A(_128_), .B(_1044_), .Y(_12_) );
XNOR2X1 XNOR2X1_16 ( .A(_12_), .B(_508_), .Y(_13_) );
INVX1 INVX1_155 ( .A(_13_), .Y(_14_) );
OR2X2 OR2X2_14 ( .A(_14_), .B(_11_), .Y(_15_) );
NAND2X1 NAND2X1_131 ( .A(_11_), .B(_14_), .Y(_16_) );
AOI21X1 AOI21X1_74 ( .A(_15_), .B(_16_), .C(_9_), .Y(_17_) );
NAND3X1 NAND3X1_117 ( .A(_9_), .B(_16_), .C(_15_), .Y(_18_) );
INVX1 INVX1_156 ( .A(_18_), .Y(_19_) );
NOR2X1 NOR2X1_151 ( .A(_17_), .B(_19_), .Y(_20_) );
XNOR2X1 XNOR2X1_17 ( .A(_20_), .B(_3_), .Y(_22_) );
XOR2X1 XOR2X1_38 ( .A(_22_), .B(_0_), .Y(_23_) );
NOR2X1 NOR2X1_152 ( .A(_1064_), .B(_23_), .Y(_24_) );
NAND2X1 NAND2X1_132 ( .A(_1064_), .B(_23_), .Y(_25_) );
INVX1 INVX1_157 ( .A(_25_), .Y(_26_) );
NOR2X1 NOR2X1_153 ( .A(_24_), .B(_26_), .Y(_27_) );
NAND2X1 NAND2X1_133 ( .A(_27_), .B(_1062_), .Y(_28_) );
INVX1 INVX1_158 ( .A(_28_), .Y(_29_) );
NOR2X1 NOR2X1_154 ( .A(_592_), .B(_29_), .Y(_30_) );
OAI21X1 OAI21X1_228 ( .A(_1062_), .B(_27_), .C(_30_), .Y(_31_) );
AOI21X1 AOI21X1_75 ( .A(_31_), .B(_1019_), .C(_406_), .Y(alu_inst_alu_out_comp_10_) );
NAND2X1 NAND2X1_134 ( .A(_3_), .B(_20_), .Y(_33_) );
OAI21X1 OAI21X1_229 ( .A(_0_), .B(_22_), .C(_33_), .Y(_34_) );
NAND2X1 NAND2X1_135 ( .A(_5_), .B(_7_), .Y(_35_) );
NAND2X1 NAND2X1_136 ( .A(_4_), .B(_8_), .Y(_36_) );
NAND2X1 NAND2X1_137 ( .A(_35_), .B(_36_), .Y(_37_) );
NAND2X1 NAND2X1_138 ( .A(_16_), .B(_18_), .Y(_38_) );
NOR2X1 NOR2X1_155 ( .A(_582_), .B(_840_), .Y(_39_) );
NOR2X1 NOR2X1_156 ( .A(_593_), .B(_818_), .Y(_40_) );
NAND2X1 NAND2X1_139 ( .A(_508_), .B(_12_), .Y(_41_) );
OAI21X1 OAI21X1_230 ( .A(_128_), .B(_1044_), .C(_41_), .Y(_43_) );
XOR2X1 XOR2X1_39 ( .A(_43_), .B(_40_), .Y(_44_) );
XOR2X1 XOR2X1_40 ( .A(_44_), .B(_39_), .Y(_45_) );
INVX1 INVX1_159 ( .A(_162_), .Y(_46_) );
NOR2X1 NOR2X1_157 ( .A(_504_), .B(_505_), .Y(_47_) );
NAND2X1 NAND2X1_140 ( .A(_47_), .B(_46_), .Y(_48_) );
OAI21X1 OAI21X1_231 ( .A(_504_), .B(_505_), .C(_162_), .Y(_49_) );
AND2X2 AND2X2_33 ( .A(_48_), .B(_49_), .Y(_50_) );
XOR2X1 XOR2X1_41 ( .A(_50_), .B(_45_), .Y(_51_) );
XOR2X1 XOR2X1_42 ( .A(_51_), .B(_38_), .Y(_52_) );
XOR2X1 XOR2X1_43 ( .A(_52_), .B(_37_), .Y(_54_) );
XOR2X1 XOR2X1_44 ( .A(_54_), .B(_34_), .Y(_55_) );
OAI21X1 OAI21X1_232 ( .A(_26_), .B(_29_), .C(_55_), .Y(_56_) );
INVX1 INVX1_160 ( .A(_55_), .Y(_57_) );
NAND3X1 NAND3X1_118 ( .A(_25_), .B(_57_), .C(_28_), .Y(_58_) );
NAND3X1 NAND3X1_119 ( .A(_591_), .B(_58_), .C(_56_), .Y(_59_) );
AOI21X1 AOI21X1_76 ( .A(_59_), .B(_1019_), .C(_406_), .Y(alu_inst_alu_out_comp_11_) );
NAND2X1 NAND2X1_141 ( .A(_34_), .B(_54_), .Y(_60_) );
NAND2X1 NAND2X1_142 ( .A(_60_), .B(_56_), .Y(_61_) );
NAND2X1 NAND2X1_143 ( .A(_38_), .B(_51_), .Y(_62_) );
NAND2X1 NAND2X1_144 ( .A(_37_), .B(_52_), .Y(_64_) );
NAND2X1 NAND2X1_145 ( .A(_62_), .B(_64_), .Y(_65_) );
NAND2X1 NAND2X1_146 ( .A(_40_), .B(_43_), .Y(_66_) );
NAND2X1 NAND2X1_147 ( .A(_39_), .B(_44_), .Y(_67_) );
NAND2X1 NAND2X1_148 ( .A(_66_), .B(_67_), .Y(_68_) );
INVX1 INVX1_161 ( .A(_68_), .Y(_69_) );
NAND2X1 NAND2X1_149 ( .A(_45_), .B(_50_), .Y(_70_) );
OAI21X1 OAI21X1_233 ( .A(_593_), .B(_504_), .C(_48_), .Y(_71_) );
OAI21X1 OAI21X1_234 ( .A(_593_), .B(_48_), .C(_71_), .Y(_72_) );
OAI21X1 OAI21X1_235 ( .A(_582_), .B(_818_), .C(_72_), .Y(_73_) );
INVX1 INVX1_162 ( .A(_72_), .Y(_75_) );
NAND3X1 NAND3X1_120 ( .A(alu_inst_data_b_in_7_), .B(alu_inst_data_a_in_5_), .C(_75_), .Y(_76_) );
AND2X2 AND2X2_34 ( .A(_76_), .B(_73_), .Y(_77_) );
INVX1 INVX1_163 ( .A(_77_), .Y(_78_) );
OR2X2 OR2X2_15 ( .A(_78_), .B(_237_), .Y(_79_) );
OAI21X1 OAI21X1_236 ( .A(_505_), .B(_224_), .C(_78_), .Y(_80_) );
NAND2X1 NAND2X1_150 ( .A(_80_), .B(_79_), .Y(_81_) );
NAND2X1 NAND2X1_151 ( .A(_70_), .B(_81_), .Y(_82_) );
OR2X2 OR2X2_16 ( .A(_81_), .B(_70_), .Y(_83_) );
NAND2X1 NAND2X1_152 ( .A(_82_), .B(_83_), .Y(_84_) );
XOR2X1 XOR2X1_45 ( .A(_84_), .B(_69_), .Y(_86_) );
NOR2X1 NOR2X1_158 ( .A(_65_), .B(_86_), .Y(_87_) );
NAND2X1 NAND2X1_153 ( .A(_65_), .B(_86_), .Y(_88_) );
INVX1 INVX1_164 ( .A(_88_), .Y(_89_) );
NOR2X1 NOR2X1_159 ( .A(_87_), .B(_89_), .Y(_90_) );
NAND2X1 NAND2X1_154 ( .A(_61_), .B(_90_), .Y(_91_) );
INVX1 INVX1_165 ( .A(_91_), .Y(_92_) );
NOR2X1 NOR2X1_160 ( .A(_592_), .B(_92_), .Y(_93_) );
OAI21X1 OAI21X1_237 ( .A(_61_), .B(_90_), .C(_93_), .Y(_94_) );
AOI21X1 AOI21X1_77 ( .A(_94_), .B(_1019_), .C(_406_), .Y(alu_inst_alu_out_comp_12_) );
OAI21X1 OAI21X1_238 ( .A(_69_), .B(_84_), .C(_83_), .Y(_96_) );
OAI21X1 OAI21X1_239 ( .A(_593_), .B(_48_), .C(_76_), .Y(_97_) );
NOR2X1 NOR2X1_161 ( .A(_582_), .B(_504_), .Y(_98_) );
NAND3X1 NAND3X1_121 ( .A(alu_inst_data_b_in_6_), .B(_98_), .C(_296_), .Y(_99_) );
INVX1 INVX1_166 ( .A(_98_), .Y(_100_) );
OAI21X1 OAI21X1_240 ( .A(_593_), .B(_297_), .C(_100_), .Y(_101_) );
NAND2X1 NAND2X1_155 ( .A(_99_), .B(_101_), .Y(_102_) );
XOR2X1 XOR2X1_46 ( .A(_102_), .B(_79_), .Y(_103_) );
OR2X2 OR2X2_17 ( .A(_103_), .B(_97_), .Y(_104_) );
NAND2X1 NAND2X1_156 ( .A(_97_), .B(_103_), .Y(_105_) );
AND2X2 AND2X2_35 ( .A(_104_), .B(_105_), .Y(_107_) );
NOR2X1 NOR2X1_162 ( .A(_96_), .B(_107_), .Y(_108_) );
NAND2X1 NAND2X1_157 ( .A(_96_), .B(_107_), .Y(_109_) );
INVX1 INVX1_167 ( .A(_109_), .Y(_110_) );
NOR2X1 NOR2X1_163 ( .A(_108_), .B(_110_), .Y(_111_) );
OAI21X1 OAI21X1_241 ( .A(_89_), .B(_92_), .C(_111_), .Y(_112_) );
NOR2X1 NOR2X1_164 ( .A(_89_), .B(_92_), .Y(_113_) );
OAI21X1 OAI21X1_242 ( .A(_108_), .B(_110_), .C(_113_), .Y(_114_) );
NAND3X1 NAND3X1_122 ( .A(_591_), .B(_114_), .C(_112_), .Y(_115_) );
AOI21X1 AOI21X1_78 ( .A(_115_), .B(_1019_), .C(_406_), .Y(alu_inst_alu_out_comp_13_) );
OAI21X1 OAI21X1_243 ( .A(_113_), .B(_108_), .C(_109_), .Y(_117_) );
OAI21X1 OAI21X1_244 ( .A(_79_), .B(_102_), .C(_105_), .Y(_118_) );
NAND2X1 NAND2X1_158 ( .A(_543_), .B(_99_), .Y(_119_) );
XNOR2X1 XNOR2X1_18 ( .A(_118_), .B(_119_), .Y(_120_) );
AOI21X1 AOI21X1_79 ( .A(_117_), .B(_120_), .C(_592_), .Y(_121_) );
OAI21X1 OAI21X1_245 ( .A(_117_), .B(_120_), .C(_121_), .Y(_122_) );
AOI21X1 AOI21X1_80 ( .A(_122_), .B(_1019_), .C(_406_), .Y(alu_inst_alu_out_comp_14_) );
AND2X2 AND2X2_36 ( .A(_117_), .B(_120_), .Y(_123_) );
NAND3X1 NAND3X1_123 ( .A(_543_), .B(_99_), .C(_118_), .Y(_124_) );
NAND2X1 NAND2X1_159 ( .A(_99_), .B(_124_), .Y(_125_) );
OAI21X1 OAI21X1_246 ( .A(_125_), .B(_123_), .C(_591_), .Y(_127_) );
AOI21X1 AOI21X1_81 ( .A(_127_), .B(_1019_), .C(_406_), .Y(alu_inst_alu_out_comp_15_) );
DFFSR DFFSR_1 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_0_), .Q(alu_inst_data_out_0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_2 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_1_), .Q(alu_inst_data_out_1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_3 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_2_), .Q(alu_inst_data_out_2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_4 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_3_), .Q(alu_inst_data_out_3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_5 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_4_), .Q(alu_inst_data_out_4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_6 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_5_), .Q(alu_inst_data_out_5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_7 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_6_), .Q(alu_inst_data_out_6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_8 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_7_), .Q(alu_inst_data_out_7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_9 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_8_), .Q(alu_inst_data_out_8_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_10 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_9_), .Q(alu_inst_data_out_9_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_11 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_10_), .Q(alu_inst_data_out_10_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_12 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_11_), .Q(alu_inst_data_out_11_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_13 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_12_), .Q(alu_inst_data_out_12_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_14 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_13_), .Q(alu_inst_data_out_13_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_15 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_14_), .Q(alu_inst_data_out_14_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_16 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_15_), .Q(alu_inst_data_out_15_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_17 ( .CLK(alu_inst_clk), .D(alu_inst_alu_out_comp_valid), .Q(alu_inst_data_valid_out), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_18 ( .CLK(ref_clk), .D(bit_synchronizer_inst_reg_file_0__0_), .Q(bit_synchronizer_inst_sync_data_out), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_19 ( .CLK(ref_clk), .D(bit_synchronizer_inst_reg_file_0__1_), .Q(bit_synchronizer_inst_reg_file_0__0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_20 ( .CLK(ref_clk), .D(bit_synchronizer_inst_async_data_in), .Q(bit_synchronizer_inst_reg_file_0__1_), .R(alu_inst_reset_n), .S(_true) );
INVX1 INVX1_168 ( .A(clk_divider_inst_div_ratio_in_3_), .Y(_1069_) );
INVX1 INVX1_169 ( .A(clk_divider_inst_count_1_), .Y(_1070_) );
INVX1 INVX1_170 ( .A(clk_divider_inst_count_3_), .Y(_1071_) );
OAI22X1 OAI22X1_5 ( .A(clk_divider_inst_div_ratio_in_2_), .B(_1070_), .C(_1071_), .D(clk_divider_inst_div_ratio_in_4_), .Y(_1072_) );
AOI21X1 AOI21X1_82 ( .A(clk_divider_inst_count_2_), .B(_1069_), .C(_1072_), .Y(_1073_) );
INVX1 INVX1_171 ( .A(clk_divider_inst_div_ratio_in_2_), .Y(_1074_) );
INVX1 INVX1_172 ( .A(clk_divider_inst_count_0_), .Y(_1075_) );
NOR2X1 NOR2X1_165 ( .A(clk_divider_inst_div_ratio_in_1_), .B(_1075_), .Y(_1076_) );
OAI21X1 OAI21X1_247 ( .A(clk_divider_inst_count_1_), .B(_1074_), .C(_1076_), .Y(_1077_) );
INVX1 INVX1_173 ( .A(clk_divider_inst_div_ratio_in_4_), .Y(_1078_) );
NOR2X1 NOR2X1_166 ( .A(clk_divider_inst_count_3_), .B(_1078_), .Y(_1079_) );
NOR2X1 NOR2X1_167 ( .A(clk_divider_inst_count_2_), .B(_1069_), .Y(_1080_) );
NOR2X1 NOR2X1_168 ( .A(_1079_), .B(_1080_), .Y(_1081_) );
NAND3X1 NAND3X1_124 ( .A(_1077_), .B(_1073_), .C(_1081_), .Y(_1082_) );
NAND2X1 NAND2X1_160 ( .A(clk_divider_inst_count_3_), .B(_1078_), .Y(_1083_) );
AOI21X1 AOI21X1_83 ( .A(_1080_), .B(_1083_), .C(_1079_), .Y(_1084_) );
INVX1 INVX1_174 ( .A(clk_divider_inst_count_4_), .Y(_1085_) );
NAND2X1 NAND2X1_161 ( .A(_1070_), .B(_1075_), .Y(_1086_) );
INVX1 INVX1_175 ( .A(clk_divider_inst_count_2_), .Y(_1087_) );
NAND2X1 NAND2X1_162 ( .A(_1071_), .B(_1087_), .Y(_1088_) );
OAI21X1 OAI21X1_248 ( .A(_1086_), .B(_1088_), .C(_1085_), .Y(_1089_) );
AOI21X1 AOI21X1_84 ( .A(_1082_), .B(_1084_), .C(_1089_), .Y(clk_divider_inst_div_clk_out) );
INVX1 INVX1_176 ( .A(_true), .Y(_1090_) );
OR2X2 OR2X2_18 ( .A(clk_divider_inst_count_0_), .B(clk_divider_inst_div_ratio_in_0_), .Y(_1091_) );
NAND2X1 NAND2X1_163 ( .A(clk_divider_inst_count_0_), .B(clk_divider_inst_div_ratio_in_0_), .Y(_1092_) );
NAND2X1 NAND2X1_164 ( .A(clk_divider_inst_count_3_), .B(clk_divider_inst_div_ratio_in_3_), .Y(_1093_) );
NAND2X1 NAND2X1_165 ( .A(_1071_), .B(_1069_), .Y(_1094_) );
AOI22X1 AOI22X1_21 ( .A(_1091_), .B(_1092_), .C(_1093_), .D(_1094_), .Y(_1095_) );
XNOR2X1 XNOR2X1_19 ( .A(clk_divider_inst_count_4_), .B(clk_divider_inst_div_ratio_in_4_), .Y(_1096_) );
XNOR2X1 XNOR2X1_20 ( .A(clk_divider_inst_count_1_), .B(clk_divider_inst_div_ratio_in_1_), .Y(_1097_) );
XNOR2X1 XNOR2X1_21 ( .A(clk_divider_inst_count_2_), .B(clk_divider_inst_div_ratio_in_2_), .Y(_1098_) );
AND2X2 AND2X2_37 ( .A(_1097_), .B(_1098_), .Y(_1099_) );
NAND3X1 NAND3X1_125 ( .A(_1095_), .B(_1096_), .C(_1099_), .Y(_1100_) );
AOI21X1 AOI21X1_85 ( .A(_1100_), .B(clk_divider_inst_count_0_), .C(_1090_), .Y(_1068__0_) );
NAND2X1 NAND2X1_166 ( .A(_1092_), .B(_1091_), .Y(_1101_) );
NAND2X1 NAND2X1_167 ( .A(_1097_), .B(_1101_), .Y(_1102_) );
XNOR2X1 XNOR2X1_22 ( .A(clk_divider_inst_count_3_), .B(clk_divider_inst_div_ratio_in_3_), .Y(_1103_) );
NAND3X1 NAND3X1_126 ( .A(_1103_), .B(_1096_), .C(_1098_), .Y(_1104_) );
OAI21X1 OAI21X1_249 ( .A(clk_divider_inst_count_1_), .B(clk_divider_inst_count_0_), .C(_true), .Y(_1105_) );
AOI21X1 AOI21X1_86 ( .A(clk_divider_inst_count_1_), .B(clk_divider_inst_count_0_), .C(_1105_), .Y(_1106_) );
OAI21X1 OAI21X1_250 ( .A(_1102_), .B(_1104_), .C(_1106_), .Y(_1107_) );
INVX1 INVX1_177 ( .A(_1107_), .Y(_1068__1_) );
NAND3X1 NAND3X1_127 ( .A(clk_divider_inst_count_1_), .B(clk_divider_inst_count_0_), .C(clk_divider_inst_count_2_), .Y(_1108_) );
OAI21X1 OAI21X1_251 ( .A(_1070_), .B(_1075_), .C(_1087_), .Y(_1109_) );
NAND2X1 NAND2X1_168 ( .A(_1108_), .B(_1109_), .Y(_1110_) );
NOR2X1 NOR2X1_169 ( .A(_1090_), .B(_1110_), .Y(_1111_) );
OAI21X1 OAI21X1_252 ( .A(_1102_), .B(_1104_), .C(_1111_), .Y(_1112_) );
INVX1 INVX1_178 ( .A(_1112_), .Y(_1068__2_) );
OAI21X1 OAI21X1_253 ( .A(_1071_), .B(_1108_), .C(_true), .Y(_1113_) );
AOI21X1 AOI21X1_87 ( .A(_1071_), .B(_1108_), .C(_1113_), .Y(_1114_) );
OAI21X1 OAI21X1_254 ( .A(_1102_), .B(_1104_), .C(_1114_), .Y(_1115_) );
INVX1 INVX1_179 ( .A(_1115_), .Y(_1068__3_) );
NOR2X1 NOR2X1_170 ( .A(_1071_), .B(_1108_), .Y(_1116_) );
XOR2X1 XOR2X1_47 ( .A(_1116_), .B(_1085_), .Y(_1117_) );
OAI21X1 OAI21X1_255 ( .A(_1102_), .B(_1104_), .C(_true), .Y(_1118_) );
NOR2X1 NOR2X1_171 ( .A(_1117_), .B(_1118_), .Y(_1068__4_) );
DFFSR DFFSR_21 ( .CLK(uart_clk), .D(_1068__0_), .Q(clk_divider_inst_count_0_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_22 ( .CLK(uart_clk), .D(_1068__1_), .Q(clk_divider_inst_count_1_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_23 ( .CLK(uart_clk), .D(_1068__2_), .Q(clk_divider_inst_count_2_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_24 ( .CLK(uart_clk), .D(_1068__3_), .Q(clk_divider_inst_count_3_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_25 ( .CLK(uart_clk), .D(_1068__4_), .Q(clk_divider_inst_count_4_), .R(clk_divider_inst_reset_n), .S(_true) );
AND2X2 AND2X2_38 ( .A(clk_gate_inst_latch_out), .B(ref_clk), .Y(alu_inst_clk) );
INVX1 INVX1_180 ( .A(data_synchronizer_inst_0_ff_1_), .Y(_1127_) );
NOR2X1 NOR2X1_172 ( .A(data_synchronizer_inst_0_ff_0_), .B(_1127_), .Y(data_synchronizer_inst_0_pulse_gen) );
OAI21X1 OAI21X1_256 ( .A(data_synchronizer_inst_0_ff_0_), .B(_1127_), .C(data_synchronizer_inst_0_sync_data_out_0_), .Y(_1128_) );
INVX1 INVX1_181 ( .A(data_synchronizer_inst_0_ff_0_), .Y(_1129_) );
NAND3X1 NAND3X1_128 ( .A(data_synchronizer_inst_0_ff_1_), .B(data_synchronizer_inst_0_unsync_data_in_0_), .C(_1129_), .Y(_1130_) );
NAND2X1 NAND2X1_169 ( .A(_1130_), .B(_1128_), .Y(_1119_) );
OAI21X1 OAI21X1_257 ( .A(data_synchronizer_inst_0_ff_0_), .B(_1127_), .C(data_synchronizer_inst_0_sync_data_out_1_), .Y(_1131_) );
NAND3X1 NAND3X1_129 ( .A(data_synchronizer_inst_0_ff_1_), .B(data_synchronizer_inst_0_unsync_data_in_1_), .C(_1129_), .Y(_1132_) );
NAND2X1 NAND2X1_170 ( .A(_1132_), .B(_1131_), .Y(_1120_) );
OAI21X1 OAI21X1_258 ( .A(data_synchronizer_inst_0_ff_0_), .B(_1127_), .C(data_synchronizer_inst_0_sync_data_out_2_), .Y(_1133_) );
NAND3X1 NAND3X1_130 ( .A(data_synchronizer_inst_0_ff_1_), .B(data_synchronizer_inst_0_unsync_data_in_2_), .C(_1129_), .Y(_1134_) );
NAND2X1 NAND2X1_171 ( .A(_1134_), .B(_1133_), .Y(_1121_) );
OAI21X1 OAI21X1_259 ( .A(data_synchronizer_inst_0_ff_0_), .B(_1127_), .C(data_synchronizer_inst_0_sync_data_out_3_), .Y(_1135_) );
NAND3X1 NAND3X1_131 ( .A(data_synchronizer_inst_0_ff_1_), .B(data_synchronizer_inst_0_unsync_data_in_3_), .C(_1129_), .Y(_1136_) );
NAND2X1 NAND2X1_172 ( .A(_1136_), .B(_1135_), .Y(_1122_) );
OAI21X1 OAI21X1_260 ( .A(data_synchronizer_inst_0_ff_0_), .B(_1127_), .C(data_synchronizer_inst_0_sync_data_out_4_), .Y(_1137_) );
NAND3X1 NAND3X1_132 ( .A(data_synchronizer_inst_0_ff_1_), .B(data_synchronizer_inst_0_unsync_data_in_4_), .C(_1129_), .Y(_1138_) );
NAND2X1 NAND2X1_173 ( .A(_1138_), .B(_1137_), .Y(_1123_) );
OAI21X1 OAI21X1_261 ( .A(data_synchronizer_inst_0_ff_0_), .B(_1127_), .C(data_synchronizer_inst_0_sync_data_out_5_), .Y(_1139_) );
NAND3X1 NAND3X1_133 ( .A(data_synchronizer_inst_0_ff_1_), .B(data_synchronizer_inst_0_unsync_data_in_5_), .C(_1129_), .Y(_1140_) );
NAND2X1 NAND2X1_174 ( .A(_1140_), .B(_1139_), .Y(_1124_) );
OAI21X1 OAI21X1_262 ( .A(data_synchronizer_inst_0_ff_0_), .B(_1127_), .C(data_synchronizer_inst_0_sync_data_out_6_), .Y(_1141_) );
NAND3X1 NAND3X1_134 ( .A(data_synchronizer_inst_0_ff_1_), .B(data_synchronizer_inst_0_unsync_data_in_6_), .C(_1129_), .Y(_1142_) );
NAND2X1 NAND2X1_175 ( .A(_1142_), .B(_1141_), .Y(_1125_) );
OAI21X1 OAI21X1_263 ( .A(data_synchronizer_inst_0_ff_0_), .B(_1127_), .C(data_synchronizer_inst_0_sync_data_out_7_), .Y(_1143_) );
NAND3X1 NAND3X1_135 ( .A(data_synchronizer_inst_0_ff_1_), .B(data_synchronizer_inst_0_unsync_data_in_7_), .C(_1129_), .Y(_1144_) );
NAND2X1 NAND2X1_176 ( .A(_1144_), .B(_1143_), .Y(_1126_) );
DFFSR DFFSR_26 ( .CLK(ref_clk), .D(_1119_), .Q(data_synchronizer_inst_0_sync_data_out_0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_27 ( .CLK(ref_clk), .D(_1120_), .Q(data_synchronizer_inst_0_sync_data_out_1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_28 ( .CLK(ref_clk), .D(_1121_), .Q(data_synchronizer_inst_0_sync_data_out_2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_29 ( .CLK(ref_clk), .D(_1122_), .Q(data_synchronizer_inst_0_sync_data_out_3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_30 ( .CLK(ref_clk), .D(_1123_), .Q(data_synchronizer_inst_0_sync_data_out_4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_31 ( .CLK(ref_clk), .D(_1124_), .Q(data_synchronizer_inst_0_sync_data_out_5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_32 ( .CLK(ref_clk), .D(_1125_), .Q(data_synchronizer_inst_0_sync_data_out_6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_33 ( .CLK(ref_clk), .D(_1126_), .Q(data_synchronizer_inst_0_sync_data_out_7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_34 ( .CLK(ref_clk), .D(data_synchronizer_inst_0_pulse_gen), .Q(data_synchronizer_inst_0_enable_pulse_out), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_35 ( .CLK(ref_clk), .D(data_synchronizer_inst_0_ff_1_), .Q(data_synchronizer_inst_0_ff_0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_36 ( .CLK(ref_clk), .D(data_synchronizer_inst_0_ff_2_), .Q(data_synchronizer_inst_0_ff_1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_37 ( .CLK(ref_clk), .D(data_synchronizer_inst_0_bus_enable_in), .Q(data_synchronizer_inst_0_ff_2_), .R(alu_inst_reset_n), .S(_true) );
INVX1 INVX1_182 ( .A(data_synchronizer_inst_1_ff_1_), .Y(_1153_) );
NOR2X1 NOR2X1_173 ( .A(data_synchronizer_inst_1_ff_0_), .B(_1153_), .Y(data_synchronizer_inst_1_pulse_gen) );
OAI21X1 OAI21X1_264 ( .A(data_synchronizer_inst_1_ff_0_), .B(_1153_), .C(data_synchronizer_inst_1_sync_data_out_0_), .Y(_1154_) );
INVX1 INVX1_183 ( .A(data_synchronizer_inst_1_ff_0_), .Y(_1155_) );
NAND3X1 NAND3X1_136 ( .A(data_synchronizer_inst_1_ff_1_), .B(data_synchronizer_inst_1_unsync_data_in_0_), .C(_1155_), .Y(_1156_) );
NAND2X1 NAND2X1_177 ( .A(_1156_), .B(_1154_), .Y(_1145_) );
OAI21X1 OAI21X1_265 ( .A(data_synchronizer_inst_1_ff_0_), .B(_1153_), .C(data_synchronizer_inst_1_sync_data_out_1_), .Y(_1157_) );
NAND3X1 NAND3X1_137 ( .A(data_synchronizer_inst_1_ff_1_), .B(data_synchronizer_inst_1_unsync_data_in_1_), .C(_1155_), .Y(_1158_) );
NAND2X1 NAND2X1_178 ( .A(_1158_), .B(_1157_), .Y(_1146_) );
OAI21X1 OAI21X1_266 ( .A(data_synchronizer_inst_1_ff_0_), .B(_1153_), .C(data_synchronizer_inst_1_sync_data_out_2_), .Y(_1159_) );
NAND3X1 NAND3X1_138 ( .A(data_synchronizer_inst_1_ff_1_), .B(data_synchronizer_inst_1_unsync_data_in_2_), .C(_1155_), .Y(_1160_) );
NAND2X1 NAND2X1_179 ( .A(_1160_), .B(_1159_), .Y(_1147_) );
OAI21X1 OAI21X1_267 ( .A(data_synchronizer_inst_1_ff_0_), .B(_1153_), .C(data_synchronizer_inst_1_sync_data_out_3_), .Y(_1161_) );
NAND3X1 NAND3X1_139 ( .A(data_synchronizer_inst_1_ff_1_), .B(data_synchronizer_inst_1_unsync_data_in_3_), .C(_1155_), .Y(_1162_) );
NAND2X1 NAND2X1_180 ( .A(_1162_), .B(_1161_), .Y(_1148_) );
OAI21X1 OAI21X1_268 ( .A(data_synchronizer_inst_1_ff_0_), .B(_1153_), .C(data_synchronizer_inst_1_sync_data_out_4_), .Y(_1163_) );
NAND3X1 NAND3X1_140 ( .A(data_synchronizer_inst_1_ff_1_), .B(data_synchronizer_inst_1_unsync_data_in_4_), .C(_1155_), .Y(_1164_) );
NAND2X1 NAND2X1_181 ( .A(_1164_), .B(_1163_), .Y(_1149_) );
OAI21X1 OAI21X1_269 ( .A(data_synchronizer_inst_1_ff_0_), .B(_1153_), .C(data_synchronizer_inst_1_sync_data_out_5_), .Y(_1165_) );
NAND3X1 NAND3X1_141 ( .A(data_synchronizer_inst_1_ff_1_), .B(data_synchronizer_inst_1_unsync_data_in_5_), .C(_1155_), .Y(_1166_) );
NAND2X1 NAND2X1_182 ( .A(_1166_), .B(_1165_), .Y(_1150_) );
OAI21X1 OAI21X1_270 ( .A(data_synchronizer_inst_1_ff_0_), .B(_1153_), .C(data_synchronizer_inst_1_sync_data_out_6_), .Y(_1167_) );
NAND3X1 NAND3X1_142 ( .A(data_synchronizer_inst_1_ff_1_), .B(data_synchronizer_inst_1_unsync_data_in_6_), .C(_1155_), .Y(_1168_) );
NAND2X1 NAND2X1_183 ( .A(_1168_), .B(_1167_), .Y(_1151_) );
OAI21X1 OAI21X1_271 ( .A(data_synchronizer_inst_1_ff_0_), .B(_1153_), .C(data_synchronizer_inst_1_sync_data_out_7_), .Y(_1169_) );
NAND3X1 NAND3X1_143 ( .A(data_synchronizer_inst_1_ff_1_), .B(data_synchronizer_inst_1_unsync_data_in_7_), .C(_1155_), .Y(_1170_) );
NAND2X1 NAND2X1_184 ( .A(_1170_), .B(_1169_), .Y(_1152_) );
DFFSR DFFSR_38 ( .CLK(clk_divider_inst_div_clk_out), .D(_1145_), .Q(data_synchronizer_inst_1_sync_data_out_0_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_39 ( .CLK(clk_divider_inst_div_clk_out), .D(_1146_), .Q(data_synchronizer_inst_1_sync_data_out_1_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_40 ( .CLK(clk_divider_inst_div_clk_out), .D(_1147_), .Q(data_synchronizer_inst_1_sync_data_out_2_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_41 ( .CLK(clk_divider_inst_div_clk_out), .D(_1148_), .Q(data_synchronizer_inst_1_sync_data_out_3_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_42 ( .CLK(clk_divider_inst_div_clk_out), .D(_1149_), .Q(data_synchronizer_inst_1_sync_data_out_4_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_43 ( .CLK(clk_divider_inst_div_clk_out), .D(_1150_), .Q(data_synchronizer_inst_1_sync_data_out_5_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_44 ( .CLK(clk_divider_inst_div_clk_out), .D(_1151_), .Q(data_synchronizer_inst_1_sync_data_out_6_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_45 ( .CLK(clk_divider_inst_div_clk_out), .D(_1152_), .Q(data_synchronizer_inst_1_sync_data_out_7_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_46 ( .CLK(clk_divider_inst_div_clk_out), .D(data_synchronizer_inst_1_pulse_gen), .Q(data_synchronizer_inst_1_enable_pulse_out), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_47 ( .CLK(clk_divider_inst_div_clk_out), .D(data_synchronizer_inst_1_ff_1_), .Q(data_synchronizer_inst_1_ff_0_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_48 ( .CLK(clk_divider_inst_div_clk_out), .D(data_synchronizer_inst_1_ff_2_), .Q(data_synchronizer_inst_1_ff_1_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_49 ( .CLK(clk_divider_inst_div_clk_out), .D(data_synchronizer_inst_1_bus_enable_in), .Q(data_synchronizer_inst_1_ff_2_), .R(clk_divider_inst_reset_n), .S(_true) );
INVX1 INVX1_184 ( .A(reg_file_inst_wr_data_in_0_), .Y(_1308_) );
INVX1 INVX1_185 ( .A(reg_file_inst_rd_en_in), .Y(_1309_) );
NAND2X1 NAND2X1_185 ( .A(reg_file_inst_wr_en_in), .B(_1309_), .Y(_1310_) );
INVX1 INVX1_186 ( .A(_1310_), .Y(_1311_) );
NAND2X1 NAND2X1_186 ( .A(reg_file_inst_addr_in_2_), .B(reg_file_inst_addr_in_3_), .Y(_1312_) );
NAND2X1 NAND2X1_187 ( .A(reg_file_inst_addr_in_0_), .B(reg_file_inst_addr_in_1_), .Y(_1313_) );
NOR2X1 NOR2X1_174 ( .A(_1312_), .B(_1313_), .Y(_1314_) );
AND2X2 AND2X2_39 ( .A(_1311_), .B(_1314_), .Y(_1315_) );
NOR2X1 NOR2X1_175 ( .A(reg_file_inst_mem_15__0_), .B(_1315_), .Y(_1316_) );
AOI21X1 AOI21X1_88 ( .A(_1308_), .B(_1315_), .C(_1316_), .Y(_1171_) );
INVX1 INVX1_187 ( .A(reg_file_inst_wr_data_in_1_), .Y(_1317_) );
NOR2X1 NOR2X1_176 ( .A(reg_file_inst_mem_15__1_), .B(_1315_), .Y(_1318_) );
AOI21X1 AOI21X1_89 ( .A(_1317_), .B(_1315_), .C(_1318_), .Y(_1172_) );
INVX1 INVX1_188 ( .A(reg_file_inst_wr_data_in_2_), .Y(_1319_) );
NOR2X1 NOR2X1_177 ( .A(reg_file_inst_mem_15__2_), .B(_1315_), .Y(_1320_) );
AOI21X1 AOI21X1_90 ( .A(_1319_), .B(_1315_), .C(_1320_), .Y(_1173_) );
INVX1 INVX1_189 ( .A(reg_file_inst_wr_data_in_3_), .Y(_1321_) );
NOR2X1 NOR2X1_178 ( .A(reg_file_inst_mem_15__3_), .B(_1315_), .Y(_1322_) );
AOI21X1 AOI21X1_91 ( .A(_1321_), .B(_1315_), .C(_1322_), .Y(_1174_) );
INVX1 INVX1_190 ( .A(reg_file_inst_wr_data_in_4_), .Y(_1323_) );
NOR2X1 NOR2X1_179 ( .A(reg_file_inst_mem_15__4_), .B(_1315_), .Y(_1324_) );
AOI21X1 AOI21X1_92 ( .A(_1323_), .B(_1315_), .C(_1324_), .Y(_1175_) );
INVX1 INVX1_191 ( .A(reg_file_inst_wr_data_in_5_), .Y(_1325_) );
NOR2X1 NOR2X1_180 ( .A(reg_file_inst_mem_15__5_), .B(_1315_), .Y(_1326_) );
AOI21X1 AOI21X1_93 ( .A(_1325_), .B(_1315_), .C(_1326_), .Y(_1176_) );
INVX1 INVX1_192 ( .A(reg_file_inst_wr_data_in_6_), .Y(_1327_) );
NOR2X1 NOR2X1_181 ( .A(reg_file_inst_mem_15__6_), .B(_1315_), .Y(_1328_) );
AOI21X1 AOI21X1_94 ( .A(_1327_), .B(_1315_), .C(_1328_), .Y(_1177_) );
INVX1 INVX1_193 ( .A(reg_file_inst_wr_data_in_7_), .Y(_1329_) );
NOR2X1 NOR2X1_182 ( .A(reg_file_inst_mem_15__7_), .B(_1315_), .Y(_1330_) );
AOI21X1 AOI21X1_95 ( .A(_1329_), .B(_1315_), .C(_1330_), .Y(_1178_) );
INVX1 INVX1_194 ( .A(reg_file_inst_rd_data_out_0_), .Y(_1331_) );
NOR2X1 NOR2X1_183 ( .A(reg_file_inst_wr_en_in), .B(_1309_), .Y(_1332_) );
INVX1 INVX1_195 ( .A(_1332_), .Y(_1333_) );
INVX1 INVX1_196 ( .A(uart_top_inst_par_en_in), .Y(_1334_) );
NOR2X1 NOR2X1_184 ( .A(reg_file_inst_addr_in_2_), .B(reg_file_inst_addr_in_3_), .Y(_1335_) );
INVX1 INVX1_197 ( .A(reg_file_inst_addr_in_0_), .Y(_1336_) );
NAND2X1 NAND2X1_188 ( .A(reg_file_inst_addr_in_1_), .B(_1336_), .Y(_1337_) );
INVX1 INVX1_198 ( .A(_1337_), .Y(_1338_) );
NAND2X1 NAND2X1_189 ( .A(_1335_), .B(_1338_), .Y(_1339_) );
OAI21X1 OAI21X1_272 ( .A(_1334_), .B(_1339_), .C(_1332_), .Y(_1340_) );
INVX1 INVX1_199 ( .A(reg_file_inst_mem_13__0_), .Y(_1341_) );
INVX1 INVX1_200 ( .A(reg_file_inst_mem_7__0_), .Y(_1342_) );
AND2X2 AND2X2_40 ( .A(reg_file_inst_addr_in_0_), .B(reg_file_inst_addr_in_1_), .Y(_1343_) );
INVX1 INVX1_201 ( .A(reg_file_inst_addr_in_3_), .Y(_1344_) );
NAND2X1 NAND2X1_190 ( .A(reg_file_inst_addr_in_2_), .B(_1344_), .Y(_1345_) );
INVX1 INVX1_202 ( .A(_1345_), .Y(_1346_) );
NAND2X1 NAND2X1_191 ( .A(_1343_), .B(_1346_), .Y(_1347_) );
NOR3X1 NOR3X1_3 ( .A(reg_file_inst_addr_in_1_), .B(_1336_), .C(_1312_), .Y(_1348_) );
INVX1 INVX1_203 ( .A(_1348_), .Y(_1349_) );
OAI22X1 OAI22X1_6 ( .A(_1342_), .B(_1347_), .C(_1341_), .D(_1349_), .Y(_1350_) );
INVX1 INVX1_204 ( .A(reg_file_inst_mem_12__0_), .Y(_1351_) );
INVX1 INVX1_205 ( .A(reg_file_inst_addr_in_2_), .Y(_1352_) );
NAND2X1 NAND2X1_192 ( .A(reg_file_inst_addr_in_3_), .B(_1352_), .Y(_1353_) );
NOR2X1 NOR2X1_185 ( .A(_1337_), .B(_1353_), .Y(_1354_) );
NAND2X1 NAND2X1_193 ( .A(reg_file_inst_mem_10__0_), .B(_1354_), .Y(_1355_) );
AND2X2 AND2X2_41 ( .A(reg_file_inst_addr_in_2_), .B(reg_file_inst_addr_in_3_), .Y(_1356_) );
NOR2X1 NOR2X1_186 ( .A(reg_file_inst_addr_in_0_), .B(reg_file_inst_addr_in_1_), .Y(_1357_) );
AND2X2 AND2X2_42 ( .A(_1356_), .B(_1357_), .Y(_1358_) );
INVX1 INVX1_206 ( .A(_1358_), .Y(_1359_) );
OAI21X1 OAI21X1_273 ( .A(_1351_), .B(_1359_), .C(_1355_), .Y(_1360_) );
NOR3X1 NOR3X1_4 ( .A(_1340_), .B(_1350_), .C(_1360_), .Y(_1361_) );
NOR3X1 NOR3X1_5 ( .A(reg_file_inst_addr_in_2_), .B(_1344_), .C(_1313_), .Y(_1362_) );
NAND2X1 NAND2X1_194 ( .A(reg_file_inst_mem_11__0_), .B(_1362_), .Y(_1363_) );
INVX1 INVX1_207 ( .A(reg_file_inst_addr_in_1_), .Y(_1364_) );
NAND2X1 NAND2X1_195 ( .A(reg_file_inst_addr_in_0_), .B(_1364_), .Y(_1365_) );
INVX1 INVX1_208 ( .A(_1365_), .Y(_1366_) );
NAND3X1 NAND3X1_144 ( .A(alu_inst_data_b_in_0_), .B(_1335_), .C(_1366_), .Y(_1367_) );
NAND3X1 NAND3X1_145 ( .A(reg_file_inst_mem_5__0_), .B(_1346_), .C(_1366_), .Y(_1368_) );
NAND3X1 NAND3X1_146 ( .A(_1367_), .B(_1363_), .C(_1368_), .Y(_1369_) );
AND2X2 AND2X2_43 ( .A(_1343_), .B(_1335_), .Y(_1370_) );
NOR2X1 NOR2X1_187 ( .A(_1337_), .B(_1345_), .Y(_1371_) );
AOI22X1 AOI22X1_22 ( .A(clk_divider_inst_div_ratio_in_0_), .B(_1370_), .C(_1371_), .D(reg_file_inst_mem_6__0_), .Y(_1372_) );
NAND3X1 NAND3X1_147 ( .A(reg_file_inst_mem_4__0_), .B(_1357_), .C(_1346_), .Y(_1373_) );
NOR2X1 NOR2X1_188 ( .A(_1365_), .B(_1353_), .Y(_1374_) );
NAND2X1 NAND2X1_196 ( .A(reg_file_inst_mem_9__0_), .B(_1374_), .Y(_1375_) );
NAND3X1 NAND3X1_148 ( .A(_1373_), .B(_1375_), .C(_1372_), .Y(_1376_) );
AND2X2 AND2X2_44 ( .A(_1335_), .B(_1357_), .Y(_1377_) );
AOI22X1 AOI22X1_23 ( .A(reg_file_inst_mem_15__0_), .B(_1314_), .C(_1377_), .D(alu_inst_data_a_in_0_), .Y(_1378_) );
INVX1 INVX1_209 ( .A(_1353_), .Y(_1379_) );
NAND3X1 NAND3X1_149 ( .A(reg_file_inst_mem_8__0_), .B(_1357_), .C(_1379_), .Y(_1380_) );
NOR2X1 NOR2X1_189 ( .A(_1312_), .B(_1337_), .Y(_1381_) );
NAND2X1 NAND2X1_197 ( .A(reg_file_inst_mem_14__0_), .B(_1381_), .Y(_1382_) );
NAND3X1 NAND3X1_150 ( .A(_1380_), .B(_1382_), .C(_1378_), .Y(_1383_) );
NOR3X1 NOR3X1_6 ( .A(_1369_), .B(_1383_), .C(_1376_), .Y(_1384_) );
AOI22X1 AOI22X1_24 ( .A(_1331_), .B(_1333_), .C(_1384_), .D(_1361_), .Y(_1179_) );
INVX1 INVX1_210 ( .A(reg_file_inst_rd_data_out_1_), .Y(_1385_) );
INVX1 INVX1_211 ( .A(uart_top_inst_par_type_in), .Y(_1386_) );
OAI21X1 OAI21X1_274 ( .A(_1386_), .B(_1339_), .C(_1332_), .Y(_1387_) );
INVX1 INVX1_212 ( .A(reg_file_inst_mem_13__1_), .Y(_1388_) );
INVX1 INVX1_213 ( .A(reg_file_inst_mem_7__1_), .Y(_1389_) );
OAI22X1 OAI22X1_7 ( .A(_1389_), .B(_1347_), .C(_1388_), .D(_1349_), .Y(_1390_) );
INVX1 INVX1_214 ( .A(reg_file_inst_mem_12__1_), .Y(_1391_) );
NAND2X1 NAND2X1_198 ( .A(reg_file_inst_mem_10__1_), .B(_1354_), .Y(_1392_) );
OAI21X1 OAI21X1_275 ( .A(_1391_), .B(_1359_), .C(_1392_), .Y(_1393_) );
NOR3X1 NOR3X1_7 ( .A(_1387_), .B(_1390_), .C(_1393_), .Y(_1394_) );
NAND2X1 NAND2X1_199 ( .A(reg_file_inst_mem_11__1_), .B(_1362_), .Y(_1395_) );
NAND3X1 NAND3X1_151 ( .A(alu_inst_data_b_in_1_), .B(_1335_), .C(_1366_), .Y(_1396_) );
NAND3X1 NAND3X1_152 ( .A(reg_file_inst_mem_5__1_), .B(_1346_), .C(_1366_), .Y(_1397_) );
NAND3X1 NAND3X1_153 ( .A(_1396_), .B(_1395_), .C(_1397_), .Y(_1398_) );
AOI22X1 AOI22X1_25 ( .A(clk_divider_inst_div_ratio_in_1_), .B(_1370_), .C(_1371_), .D(reg_file_inst_mem_6__1_), .Y(_1399_) );
NAND3X1 NAND3X1_154 ( .A(reg_file_inst_mem_4__1_), .B(_1357_), .C(_1346_), .Y(_1400_) );
NAND2X1 NAND2X1_200 ( .A(reg_file_inst_mem_9__1_), .B(_1374_), .Y(_1401_) );
NAND3X1 NAND3X1_155 ( .A(_1400_), .B(_1401_), .C(_1399_), .Y(_1402_) );
AOI22X1 AOI22X1_26 ( .A(reg_file_inst_mem_15__1_), .B(_1314_), .C(_1377_), .D(alu_inst_data_a_in_1_), .Y(_1403_) );
NAND3X1 NAND3X1_156 ( .A(reg_file_inst_mem_8__1_), .B(_1357_), .C(_1379_), .Y(_1404_) );
NAND2X1 NAND2X1_201 ( .A(reg_file_inst_mem_14__1_), .B(_1381_), .Y(_1405_) );
NAND3X1 NAND3X1_157 ( .A(_1404_), .B(_1405_), .C(_1403_), .Y(_1406_) );
NOR3X1 NOR3X1_8 ( .A(_1398_), .B(_1406_), .C(_1402_), .Y(_1407_) );
AOI22X1 AOI22X1_27 ( .A(_1385_), .B(_1333_), .C(_1407_), .D(_1394_), .Y(_1180_) );
INVX1 INVX1_215 ( .A(reg_file_inst_rd_data_out_2_), .Y(_1408_) );
INVX1 INVX1_216 ( .A(reg_file_inst_mem_14__2_), .Y(_1409_) );
NAND2X1 NAND2X1_202 ( .A(_1356_), .B(_1338_), .Y(_1410_) );
OAI21X1 OAI21X1_276 ( .A(_1409_), .B(_1410_), .C(_1332_), .Y(_1411_) );
INVX1 INVX1_217 ( .A(clk_divider_inst_div_ratio_in_2_), .Y(_1412_) );
INVX1 INVX1_218 ( .A(_1370_), .Y(_1413_) );
NAND2X1 NAND2X1_203 ( .A(reg_file_inst_mem_10__2_), .B(_1354_), .Y(_1414_) );
OAI21X1 OAI21X1_277 ( .A(_1412_), .B(_1413_), .C(_1414_), .Y(_1415_) );
INVX1 INVX1_219 ( .A(reg_file_inst_mem_9__2_), .Y(_1416_) );
INVX1 INVX1_220 ( .A(_1374_), .Y(_1417_) );
NAND2X1 NAND2X1_204 ( .A(reg_file_inst_mem_6__2_), .B(_1371_), .Y(_1418_) );
OAI21X1 OAI21X1_278 ( .A(_1416_), .B(_1417_), .C(_1418_), .Y(_1419_) );
NOR3X1 NOR3X1_9 ( .A(_1411_), .B(_1415_), .C(_1419_), .Y(_1420_) );
NAND3X1 NAND3X1_158 ( .A(reg_file_inst_mem_7__2_), .B(_1343_), .C(_1346_), .Y(_1421_) );
NAND3X1 NAND3X1_159 ( .A(alu_inst_data_b_in_2_), .B(_1335_), .C(_1366_), .Y(_1422_) );
NAND2X1 NAND2X1_205 ( .A(reg_file_inst_mem_11__2_), .B(_1362_), .Y(_1423_) );
NAND3X1 NAND3X1_160 ( .A(_1421_), .B(_1422_), .C(_1423_), .Y(_1424_) );
AOI22X1 AOI22X1_28 ( .A(_1348_), .B(reg_file_inst_mem_13__2_), .C(reg_file_inst_mem_12__2_), .D(_1358_), .Y(_1425_) );
NAND2X1 NAND2X1_206 ( .A(alu_inst_data_a_in_2_), .B(_1377_), .Y(_1426_) );
NAND3X1 NAND3X1_161 ( .A(reg_file_inst_mem_4__2_), .B(_1357_), .C(_1346_), .Y(_1427_) );
NAND3X1 NAND3X1_162 ( .A(_1426_), .B(_1427_), .C(_1425_), .Y(_1428_) );
OR2X2 OR2X2_19 ( .A(reg_file_inst_addr_in_0_), .B(reg_file_inst_addr_in_1_), .Y(_1429_) );
NOR2X1 NOR2X1_190 ( .A(_1429_), .B(_1353_), .Y(_1430_) );
AOI22X1 AOI22X1_29 ( .A(reg_file_inst_mem_15__2_), .B(_1314_), .C(_1430_), .D(reg_file_inst_mem_8__2_), .Y(_1431_) );
NAND3X1 NAND3X1_163 ( .A(reg_file_inst_mem_2__2_), .B(_1335_), .C(_1338_), .Y(_1432_) );
NOR2X1 NOR2X1_191 ( .A(_1345_), .B(_1365_), .Y(_1433_) );
NAND2X1 NAND2X1_207 ( .A(reg_file_inst_mem_5__2_), .B(_1433_), .Y(_1434_) );
NAND3X1 NAND3X1_164 ( .A(_1432_), .B(_1434_), .C(_1431_), .Y(_1435_) );
NOR3X1 NOR3X1_10 ( .A(_1424_), .B(_1428_), .C(_1435_), .Y(_1436_) );
AOI22X1 AOI22X1_30 ( .A(_1408_), .B(_1333_), .C(_1436_), .D(_1420_), .Y(_1181_) );
INVX1 INVX1_221 ( .A(reg_file_inst_rd_data_out_3_), .Y(_1437_) );
INVX1 INVX1_222 ( .A(reg_file_inst_mem_14__3_), .Y(_1438_) );
OAI21X1 OAI21X1_279 ( .A(_1438_), .B(_1410_), .C(_1332_), .Y(_1439_) );
INVX1 INVX1_223 ( .A(clk_divider_inst_div_ratio_in_3_), .Y(_1440_) );
NAND2X1 NAND2X1_208 ( .A(reg_file_inst_mem_10__3_), .B(_1354_), .Y(_1441_) );
OAI21X1 OAI21X1_280 ( .A(_1440_), .B(_1413_), .C(_1441_), .Y(_1442_) );
INVX1 INVX1_224 ( .A(reg_file_inst_mem_9__3_), .Y(_1443_) );
NAND2X1 NAND2X1_209 ( .A(reg_file_inst_mem_6__3_), .B(_1371_), .Y(_1444_) );
OAI21X1 OAI21X1_281 ( .A(_1443_), .B(_1417_), .C(_1444_), .Y(_1445_) );
NOR3X1 NOR3X1_11 ( .A(_1439_), .B(_1442_), .C(_1445_), .Y(_1446_) );
NAND3X1 NAND3X1_165 ( .A(reg_file_inst_mem_7__3_), .B(_1343_), .C(_1346_), .Y(_1447_) );
NAND3X1 NAND3X1_166 ( .A(alu_inst_data_b_in_3_), .B(_1335_), .C(_1366_), .Y(_1448_) );
NAND2X1 NAND2X1_210 ( .A(reg_file_inst_mem_11__3_), .B(_1362_), .Y(_1449_) );
NAND3X1 NAND3X1_167 ( .A(_1447_), .B(_1448_), .C(_1449_), .Y(_1450_) );
AOI22X1 AOI22X1_31 ( .A(_1348_), .B(reg_file_inst_mem_13__3_), .C(reg_file_inst_mem_12__3_), .D(_1358_), .Y(_1451_) );
NAND2X1 NAND2X1_211 ( .A(alu_inst_data_a_in_3_), .B(_1377_), .Y(_1452_) );
NAND3X1 NAND3X1_168 ( .A(reg_file_inst_mem_4__3_), .B(_1357_), .C(_1346_), .Y(_1453_) );
NAND3X1 NAND3X1_169 ( .A(_1452_), .B(_1453_), .C(_1451_), .Y(_1454_) );
AOI22X1 AOI22X1_32 ( .A(reg_file_inst_mem_15__3_), .B(_1314_), .C(_1430_), .D(reg_file_inst_mem_8__3_), .Y(_1455_) );
NAND3X1 NAND3X1_170 ( .A(reg_file_inst_mem_2__3_), .B(_1335_), .C(_1338_), .Y(_1456_) );
NAND2X1 NAND2X1_212 ( .A(reg_file_inst_mem_5__3_), .B(_1433_), .Y(_1457_) );
NAND3X1 NAND3X1_171 ( .A(_1456_), .B(_1457_), .C(_1455_), .Y(_1458_) );
NOR3X1 NOR3X1_12 ( .A(_1450_), .B(_1454_), .C(_1458_), .Y(_1459_) );
AOI22X1 AOI22X1_33 ( .A(_1437_), .B(_1333_), .C(_1459_), .D(_1446_), .Y(_1182_) );
INVX1 INVX1_225 ( .A(reg_file_inst_rd_data_out_4_), .Y(_1460_) );
INVX1 INVX1_226 ( .A(reg_file_inst_mem_2__4_), .Y(_1461_) );
OAI21X1 OAI21X1_282 ( .A(_1461_), .B(_1339_), .C(_1332_), .Y(_1462_) );
INVX1 INVX1_227 ( .A(reg_file_inst_mem_13__4_), .Y(_1463_) );
INVX1 INVX1_228 ( .A(reg_file_inst_mem_7__4_), .Y(_1464_) );
OAI22X1 OAI22X1_8 ( .A(_1464_), .B(_1347_), .C(_1463_), .D(_1349_), .Y(_1465_) );
INVX1 INVX1_229 ( .A(reg_file_inst_mem_12__4_), .Y(_1466_) );
NAND2X1 NAND2X1_213 ( .A(reg_file_inst_mem_10__4_), .B(_1354_), .Y(_1467_) );
OAI21X1 OAI21X1_283 ( .A(_1466_), .B(_1359_), .C(_1467_), .Y(_1468_) );
NOR3X1 NOR3X1_13 ( .A(_1462_), .B(_1465_), .C(_1468_), .Y(_1469_) );
NAND3X1 NAND3X1_172 ( .A(reg_file_inst_mem_8__4_), .B(_1357_), .C(_1379_), .Y(_1470_) );
NAND3X1 NAND3X1_173 ( .A(alu_inst_data_b_in_4_), .B(_1335_), .C(_1366_), .Y(_1471_) );
NAND3X1 NAND3X1_174 ( .A(reg_file_inst_mem_5__4_), .B(_1346_), .C(_1366_), .Y(_1472_) );
NAND3X1 NAND3X1_175 ( .A(_1470_), .B(_1471_), .C(_1472_), .Y(_1473_) );
AOI22X1 AOI22X1_34 ( .A(clk_divider_inst_div_ratio_in_4_), .B(_1370_), .C(_1371_), .D(reg_file_inst_mem_6__4_), .Y(_1474_) );
NAND3X1 NAND3X1_176 ( .A(reg_file_inst_mem_4__4_), .B(_1357_), .C(_1346_), .Y(_1475_) );
NAND2X1 NAND2X1_214 ( .A(reg_file_inst_mem_9__4_), .B(_1374_), .Y(_1476_) );
NAND3X1 NAND3X1_177 ( .A(_1475_), .B(_1476_), .C(_1474_), .Y(_1477_) );
AOI22X1 AOI22X1_35 ( .A(reg_file_inst_mem_15__4_), .B(_1314_), .C(_1377_), .D(alu_inst_data_a_in_4_), .Y(_1478_) );
NAND2X1 NAND2X1_215 ( .A(reg_file_inst_mem_11__4_), .B(_1362_), .Y(_1479_) );
NAND2X1 NAND2X1_216 ( .A(reg_file_inst_mem_14__4_), .B(_1381_), .Y(_1480_) );
NAND3X1 NAND3X1_178 ( .A(_1479_), .B(_1480_), .C(_1478_), .Y(_1481_) );
NOR3X1 NOR3X1_14 ( .A(_1473_), .B(_1481_), .C(_1477_), .Y(_1482_) );
AOI22X1 AOI22X1_36 ( .A(_1460_), .B(_1333_), .C(_1482_), .D(_1469_), .Y(_1183_) );
INVX1 INVX1_230 ( .A(reg_file_inst_rd_data_out_5_), .Y(_1483_) );
INVX1 INVX1_231 ( .A(reg_file_inst_mem_14__5_), .Y(_1484_) );
OAI21X1 OAI21X1_284 ( .A(_1484_), .B(_1410_), .C(_1332_), .Y(_1485_) );
INVX1 INVX1_232 ( .A(reg_file_inst_mem_3__5_), .Y(_1486_) );
NAND2X1 NAND2X1_217 ( .A(reg_file_inst_mem_10__5_), .B(_1354_), .Y(_1487_) );
OAI21X1 OAI21X1_285 ( .A(_1486_), .B(_1413_), .C(_1487_), .Y(_1488_) );
INVX1 INVX1_233 ( .A(reg_file_inst_mem_9__5_), .Y(_1489_) );
NAND2X1 NAND2X1_218 ( .A(reg_file_inst_mem_6__5_), .B(_1371_), .Y(_1490_) );
OAI21X1 OAI21X1_286 ( .A(_1489_), .B(_1417_), .C(_1490_), .Y(_1491_) );
NOR3X1 NOR3X1_15 ( .A(_1485_), .B(_1488_), .C(_1491_), .Y(_1492_) );
NAND3X1 NAND3X1_179 ( .A(reg_file_inst_mem_7__5_), .B(_1343_), .C(_1346_), .Y(_1493_) );
NAND3X1 NAND3X1_180 ( .A(alu_inst_data_b_in_5_), .B(_1335_), .C(_1366_), .Y(_1494_) );
NAND3X1 NAND3X1_181 ( .A(reg_file_inst_mem_8__5_), .B(_1357_), .C(_1379_), .Y(_1495_) );
NAND3X1 NAND3X1_182 ( .A(_1493_), .B(_1494_), .C(_1495_), .Y(_1496_) );
AOI22X1 AOI22X1_37 ( .A(_1348_), .B(reg_file_inst_mem_13__5_), .C(reg_file_inst_mem_12__5_), .D(_1358_), .Y(_1497_) );
NAND2X1 NAND2X1_219 ( .A(alu_inst_data_a_in_5_), .B(_1377_), .Y(_1498_) );
NAND3X1 NAND3X1_183 ( .A(reg_file_inst_mem_4__5_), .B(_1357_), .C(_1346_), .Y(_1499_) );
NAND3X1 NAND3X1_184 ( .A(_1498_), .B(_1499_), .C(_1497_), .Y(_1500_) );
AOI22X1 AOI22X1_38 ( .A(reg_file_inst_mem_15__5_), .B(_1314_), .C(_1362_), .D(reg_file_inst_mem_11__5_), .Y(_1501_) );
NAND3X1 NAND3X1_185 ( .A(reg_file_inst_mem_2__5_), .B(_1335_), .C(_1338_), .Y(_1502_) );
NAND2X1 NAND2X1_220 ( .A(reg_file_inst_mem_5__5_), .B(_1433_), .Y(_1503_) );
NAND3X1 NAND3X1_186 ( .A(_1502_), .B(_1501_), .C(_1503_), .Y(_1504_) );
NOR3X1 NOR3X1_16 ( .A(_1496_), .B(_1504_), .C(_1500_), .Y(_1505_) );
AOI22X1 AOI22X1_39 ( .A(_1483_), .B(_1333_), .C(_1505_), .D(_1492_), .Y(_1184_) );
INVX1 INVX1_234 ( .A(reg_file_inst_rd_data_out_6_), .Y(_1506_) );
INVX1 INVX1_235 ( .A(reg_file_inst_mem_14__6_), .Y(_1507_) );
OAI21X1 OAI21X1_287 ( .A(_1507_), .B(_1410_), .C(_1332_), .Y(_1508_) );
INVX1 INVX1_236 ( .A(reg_file_inst_mem_3__6_), .Y(_1509_) );
NAND2X1 NAND2X1_221 ( .A(reg_file_inst_mem_10__6_), .B(_1354_), .Y(_1510_) );
OAI21X1 OAI21X1_288 ( .A(_1509_), .B(_1413_), .C(_1510_), .Y(_1511_) );
INVX1 INVX1_237 ( .A(reg_file_inst_mem_9__6_), .Y(_1512_) );
NAND2X1 NAND2X1_222 ( .A(reg_file_inst_mem_6__6_), .B(_1371_), .Y(_1513_) );
OAI21X1 OAI21X1_289 ( .A(_1512_), .B(_1417_), .C(_1513_), .Y(_1514_) );
NOR3X1 NOR3X1_17 ( .A(_1508_), .B(_1511_), .C(_1514_), .Y(_1515_) );
NAND3X1 NAND3X1_187 ( .A(reg_file_inst_mem_7__6_), .B(_1343_), .C(_1346_), .Y(_1516_) );
NAND3X1 NAND3X1_188 ( .A(alu_inst_data_b_in_6_), .B(_1335_), .C(_1366_), .Y(_1517_) );
NAND2X1 NAND2X1_223 ( .A(reg_file_inst_mem_11__6_), .B(_1362_), .Y(_1518_) );
NAND3X1 NAND3X1_189 ( .A(_1516_), .B(_1517_), .C(_1518_), .Y(_1519_) );
AOI22X1 AOI22X1_40 ( .A(_1348_), .B(reg_file_inst_mem_13__6_), .C(reg_file_inst_mem_12__6_), .D(_1358_), .Y(_1520_) );
NAND2X1 NAND2X1_224 ( .A(alu_inst_data_a_in_6_), .B(_1377_), .Y(_1521_) );
NAND3X1 NAND3X1_190 ( .A(reg_file_inst_mem_4__6_), .B(_1357_), .C(_1346_), .Y(_1522_) );
NAND3X1 NAND3X1_191 ( .A(_1521_), .B(_1522_), .C(_1520_), .Y(_1523_) );
AOI22X1 AOI22X1_41 ( .A(reg_file_inst_mem_15__6_), .B(_1314_), .C(_1430_), .D(reg_file_inst_mem_8__6_), .Y(_1524_) );
NAND3X1 NAND3X1_192 ( .A(reg_file_inst_mem_2__6_), .B(_1335_), .C(_1338_), .Y(_1525_) );
NAND2X1 NAND2X1_225 ( .A(reg_file_inst_mem_5__6_), .B(_1433_), .Y(_1526_) );
NAND3X1 NAND3X1_193 ( .A(_1525_), .B(_1526_), .C(_1524_), .Y(_1527_) );
NOR3X1 NOR3X1_18 ( .A(_1519_), .B(_1523_), .C(_1527_), .Y(_1528_) );
AOI22X1 AOI22X1_42 ( .A(_1506_), .B(_1333_), .C(_1528_), .D(_1515_), .Y(_1185_) );
INVX1 INVX1_238 ( .A(reg_file_inst_rd_data_out_7_), .Y(_1529_) );
INVX1 INVX1_239 ( .A(reg_file_inst_mem_2__7_), .Y(_1530_) );
OAI21X1 OAI21X1_290 ( .A(_1530_), .B(_1339_), .C(_1332_), .Y(_1531_) );
INVX1 INVX1_240 ( .A(reg_file_inst_mem_13__7_), .Y(_1532_) );
INVX1 INVX1_241 ( .A(reg_file_inst_mem_7__7_), .Y(_1533_) );
OAI22X1 OAI22X1_9 ( .A(_1533_), .B(_1347_), .C(_1532_), .D(_1349_), .Y(_1534_) );
INVX1 INVX1_242 ( .A(reg_file_inst_mem_12__7_), .Y(_1535_) );
NAND2X1 NAND2X1_226 ( .A(reg_file_inst_mem_10__7_), .B(_1354_), .Y(_1536_) );
OAI21X1 OAI21X1_291 ( .A(_1535_), .B(_1359_), .C(_1536_), .Y(_1537_) );
NOR3X1 NOR3X1_19 ( .A(_1531_), .B(_1534_), .C(_1537_), .Y(_1538_) );
NAND2X1 NAND2X1_227 ( .A(reg_file_inst_mem_11__7_), .B(_1362_), .Y(_1539_) );
NAND3X1 NAND3X1_194 ( .A(alu_inst_data_b_in_7_), .B(_1335_), .C(_1366_), .Y(_1540_) );
NAND3X1 NAND3X1_195 ( .A(reg_file_inst_mem_5__7_), .B(_1346_), .C(_1366_), .Y(_1541_) );
NAND3X1 NAND3X1_196 ( .A(_1540_), .B(_1539_), .C(_1541_), .Y(_1542_) );
AOI22X1 AOI22X1_43 ( .A(reg_file_inst_mem_3__7_), .B(_1370_), .C(_1371_), .D(reg_file_inst_mem_6__7_), .Y(_1543_) );
NAND3X1 NAND3X1_197 ( .A(reg_file_inst_mem_4__7_), .B(_1357_), .C(_1346_), .Y(_1544_) );
NAND2X1 NAND2X1_228 ( .A(reg_file_inst_mem_9__7_), .B(_1374_), .Y(_1545_) );
NAND3X1 NAND3X1_198 ( .A(_1544_), .B(_1545_), .C(_1543_), .Y(_1546_) );
AOI22X1 AOI22X1_44 ( .A(reg_file_inst_mem_15__7_), .B(_1314_), .C(_1377_), .D(alu_inst_data_a_in_7_), .Y(_1547_) );
NAND3X1 NAND3X1_199 ( .A(reg_file_inst_mem_8__7_), .B(_1357_), .C(_1379_), .Y(_1548_) );
NAND2X1 NAND2X1_229 ( .A(reg_file_inst_mem_14__7_), .B(_1381_), .Y(_1549_) );
NAND3X1 NAND3X1_200 ( .A(_1548_), .B(_1549_), .C(_1547_), .Y(_1550_) );
NOR3X1 NOR3X1_20 ( .A(_1542_), .B(_1550_), .C(_1546_), .Y(_1551_) );
AOI22X1 AOI22X1_45 ( .A(_1529_), .B(_1333_), .C(_1551_), .D(_1538_), .Y(_1186_) );
AND2X2 AND2X2_45 ( .A(_1377_), .B(_1311_), .Y(_1552_) );
NOR2X1 NOR2X1_192 ( .A(alu_inst_data_a_in_0_), .B(_1552_), .Y(_1553_) );
AOI21X1 AOI21X1_96 ( .A(_1308_), .B(_1552_), .C(_1553_), .Y(_1188_) );
NOR2X1 NOR2X1_193 ( .A(alu_inst_data_a_in_1_), .B(_1552_), .Y(_1554_) );
AOI21X1 AOI21X1_97 ( .A(_1317_), .B(_1552_), .C(_1554_), .Y(_1189_) );
NOR2X1 NOR2X1_194 ( .A(alu_inst_data_a_in_2_), .B(_1552_), .Y(_1555_) );
AOI21X1 AOI21X1_98 ( .A(_1319_), .B(_1552_), .C(_1555_), .Y(_1190_) );
NOR2X1 NOR2X1_195 ( .A(alu_inst_data_a_in_3_), .B(_1552_), .Y(_1556_) );
AOI21X1 AOI21X1_99 ( .A(_1321_), .B(_1552_), .C(_1556_), .Y(_1191_) );
NOR2X1 NOR2X1_196 ( .A(alu_inst_data_a_in_4_), .B(_1552_), .Y(_1557_) );
AOI21X1 AOI21X1_100 ( .A(_1323_), .B(_1552_), .C(_1557_), .Y(_1192_) );
NOR2X1 NOR2X1_197 ( .A(alu_inst_data_a_in_5_), .B(_1552_), .Y(_1558_) );
AOI21X1 AOI21X1_101 ( .A(_1325_), .B(_1552_), .C(_1558_), .Y(_1193_) );
NOR2X1 NOR2X1_198 ( .A(alu_inst_data_a_in_6_), .B(_1552_), .Y(_1559_) );
AOI21X1 AOI21X1_102 ( .A(_1327_), .B(_1552_), .C(_1559_), .Y(_1194_) );
NOR2X1 NOR2X1_199 ( .A(alu_inst_data_a_in_7_), .B(_1552_), .Y(_1560_) );
AOI21X1 AOI21X1_103 ( .A(_1329_), .B(_1552_), .C(_1560_), .Y(_1195_) );
NAND3X1 NAND3X1_201 ( .A(_1335_), .B(_1366_), .C(_1311_), .Y(_1561_) );
NAND2X1 NAND2X1_230 ( .A(alu_inst_data_b_in_0_), .B(_1561_), .Y(_1562_) );
OAI21X1 OAI21X1_292 ( .A(_1308_), .B(_1561_), .C(_1562_), .Y(_1196_) );
NAND2X1 NAND2X1_231 ( .A(alu_inst_data_b_in_1_), .B(_1561_), .Y(_1563_) );
OAI21X1 OAI21X1_293 ( .A(_1317_), .B(_1561_), .C(_1563_), .Y(_1197_) );
NAND2X1 NAND2X1_232 ( .A(alu_inst_data_b_in_2_), .B(_1561_), .Y(_1564_) );
OAI21X1 OAI21X1_294 ( .A(_1319_), .B(_1561_), .C(_1564_), .Y(_1198_) );
NAND2X1 NAND2X1_233 ( .A(alu_inst_data_b_in_3_), .B(_1561_), .Y(_1565_) );
OAI21X1 OAI21X1_295 ( .A(_1321_), .B(_1561_), .C(_1565_), .Y(_1199_) );
NAND2X1 NAND2X1_234 ( .A(alu_inst_data_b_in_4_), .B(_1561_), .Y(_1566_) );
OAI21X1 OAI21X1_296 ( .A(_1323_), .B(_1561_), .C(_1566_), .Y(_1200_) );
NAND2X1 NAND2X1_235 ( .A(alu_inst_data_b_in_5_), .B(_1561_), .Y(_1567_) );
OAI21X1 OAI21X1_297 ( .A(_1325_), .B(_1561_), .C(_1567_), .Y(_1201_) );
NAND2X1 NAND2X1_236 ( .A(alu_inst_data_b_in_6_), .B(_1561_), .Y(_1568_) );
OAI21X1 OAI21X1_298 ( .A(_1327_), .B(_1561_), .C(_1568_), .Y(_1202_) );
NAND2X1 NAND2X1_237 ( .A(alu_inst_data_b_in_7_), .B(_1561_), .Y(_1569_) );
OAI21X1 OAI21X1_299 ( .A(_1329_), .B(_1561_), .C(_1569_), .Y(_1203_) );
NOR2X1 NOR2X1_200 ( .A(_1310_), .B(_1339_), .Y(_1570_) );
NAND2X1 NAND2X1_238 ( .A(reg_file_inst_wr_data_in_0_), .B(_1570_), .Y(_1571_) );
OAI21X1 OAI21X1_300 ( .A(_1334_), .B(_1570_), .C(_1571_), .Y(_1204_) );
NAND2X1 NAND2X1_239 ( .A(reg_file_inst_wr_data_in_1_), .B(_1570_), .Y(_1572_) );
OAI21X1 OAI21X1_301 ( .A(_1386_), .B(_1570_), .C(_1572_), .Y(_1205_) );
NOR2X1 NOR2X1_201 ( .A(reg_file_inst_mem_2__2_), .B(_1570_), .Y(_1573_) );
AOI21X1 AOI21X1_104 ( .A(_1319_), .B(_1570_), .C(_1573_), .Y(_1206_) );
NOR2X1 NOR2X1_202 ( .A(reg_file_inst_mem_2__3_), .B(_1570_), .Y(_1574_) );
AOI21X1 AOI21X1_105 ( .A(_1321_), .B(_1570_), .C(_1574_), .Y(_1207_) );
NAND2X1 NAND2X1_240 ( .A(reg_file_inst_wr_data_in_4_), .B(_1570_), .Y(_1575_) );
OAI21X1 OAI21X1_302 ( .A(_1461_), .B(_1570_), .C(_1575_), .Y(_1208_) );
NOR2X1 NOR2X1_203 ( .A(reg_file_inst_mem_2__5_), .B(_1570_), .Y(_1576_) );
AOI21X1 AOI21X1_106 ( .A(_1325_), .B(_1570_), .C(_1576_), .Y(_1209_) );
NOR2X1 NOR2X1_204 ( .A(reg_file_inst_mem_2__6_), .B(_1570_), .Y(_1577_) );
AOI21X1 AOI21X1_107 ( .A(_1327_), .B(_1570_), .C(_1577_), .Y(_1210_) );
NAND2X1 NAND2X1_241 ( .A(reg_file_inst_wr_data_in_7_), .B(_1570_), .Y(_1578_) );
OAI21X1 OAI21X1_303 ( .A(_1530_), .B(_1570_), .C(_1578_), .Y(_1211_) );
NAND2X1 NAND2X1_242 ( .A(_1311_), .B(_1370_), .Y(_1579_) );
OAI21X1 OAI21X1_304 ( .A(_1310_), .B(_1413_), .C(clk_divider_inst_div_ratio_in_0_), .Y(_1580_) );
OAI21X1 OAI21X1_305 ( .A(_1308_), .B(_1579_), .C(_1580_), .Y(_1212_) );
OAI21X1 OAI21X1_306 ( .A(_1310_), .B(_1413_), .C(clk_divider_inst_div_ratio_in_1_), .Y(_1581_) );
OAI21X1 OAI21X1_307 ( .A(_1317_), .B(_1579_), .C(_1581_), .Y(_1213_) );
OAI21X1 OAI21X1_308 ( .A(_1310_), .B(_1413_), .C(clk_divider_inst_div_ratio_in_2_), .Y(_1582_) );
OAI21X1 OAI21X1_309 ( .A(_1319_), .B(_1579_), .C(_1582_), .Y(_1214_) );
OAI21X1 OAI21X1_310 ( .A(_1310_), .B(_1413_), .C(clk_divider_inst_div_ratio_in_3_), .Y(_1583_) );
OAI21X1 OAI21X1_311 ( .A(_1321_), .B(_1579_), .C(_1583_), .Y(_1215_) );
OAI21X1 OAI21X1_312 ( .A(_1310_), .B(_1413_), .C(clk_divider_inst_div_ratio_in_4_), .Y(_1584_) );
OAI21X1 OAI21X1_313 ( .A(_1323_), .B(_1579_), .C(_1584_), .Y(_1216_) );
OAI21X1 OAI21X1_314 ( .A(_1310_), .B(_1413_), .C(reg_file_inst_mem_3__5_), .Y(_1585_) );
OAI21X1 OAI21X1_315 ( .A(_1325_), .B(_1579_), .C(_1585_), .Y(_1217_) );
OAI21X1 OAI21X1_316 ( .A(_1310_), .B(_1413_), .C(reg_file_inst_mem_3__6_), .Y(_1586_) );
OAI21X1 OAI21X1_317 ( .A(_1327_), .B(_1579_), .C(_1586_), .Y(_1218_) );
OAI21X1 OAI21X1_318 ( .A(_1310_), .B(_1413_), .C(reg_file_inst_mem_3__7_), .Y(_1587_) );
OAI21X1 OAI21X1_319 ( .A(_1329_), .B(_1579_), .C(_1587_), .Y(_1219_) );
NAND2X1 NAND2X1_243 ( .A(_1357_), .B(_1346_), .Y(_1588_) );
NOR2X1 NOR2X1_205 ( .A(_1310_), .B(_1588_), .Y(_1589_) );
NOR2X1 NOR2X1_206 ( .A(reg_file_inst_mem_4__0_), .B(_1589_), .Y(_1590_) );
AOI21X1 AOI21X1_108 ( .A(_1308_), .B(_1589_), .C(_1590_), .Y(_1220_) );
NOR2X1 NOR2X1_207 ( .A(reg_file_inst_mem_4__1_), .B(_1589_), .Y(_1591_) );
AOI21X1 AOI21X1_109 ( .A(_1317_), .B(_1589_), .C(_1591_), .Y(_1221_) );
NOR2X1 NOR2X1_208 ( .A(reg_file_inst_mem_4__2_), .B(_1589_), .Y(_1592_) );
AOI21X1 AOI21X1_110 ( .A(_1319_), .B(_1589_), .C(_1592_), .Y(_1222_) );
NOR2X1 NOR2X1_209 ( .A(reg_file_inst_mem_4__3_), .B(_1589_), .Y(_1593_) );
AOI21X1 AOI21X1_111 ( .A(_1321_), .B(_1589_), .C(_1593_), .Y(_1223_) );
NOR2X1 NOR2X1_210 ( .A(reg_file_inst_mem_4__4_), .B(_1589_), .Y(_1594_) );
AOI21X1 AOI21X1_112 ( .A(_1323_), .B(_1589_), .C(_1594_), .Y(_1224_) );
NOR2X1 NOR2X1_211 ( .A(reg_file_inst_mem_4__5_), .B(_1589_), .Y(_1595_) );
AOI21X1 AOI21X1_113 ( .A(_1325_), .B(_1589_), .C(_1595_), .Y(_1225_) );
NOR2X1 NOR2X1_212 ( .A(reg_file_inst_mem_4__6_), .B(_1589_), .Y(_1596_) );
AOI21X1 AOI21X1_114 ( .A(_1327_), .B(_1589_), .C(_1596_), .Y(_1226_) );
NOR2X1 NOR2X1_213 ( .A(reg_file_inst_mem_4__7_), .B(_1589_), .Y(_1597_) );
AOI21X1 AOI21X1_115 ( .A(_1329_), .B(_1589_), .C(_1597_), .Y(_1227_) );
NAND2X1 NAND2X1_244 ( .A(_1311_), .B(_1433_), .Y(_1598_) );
NAND2X1 NAND2X1_245 ( .A(reg_file_inst_mem_5__0_), .B(_1598_), .Y(_1599_) );
OAI21X1 OAI21X1_320 ( .A(_1308_), .B(_1598_), .C(_1599_), .Y(_1228_) );
NAND2X1 NAND2X1_246 ( .A(reg_file_inst_mem_5__1_), .B(_1598_), .Y(_1600_) );
OAI21X1 OAI21X1_321 ( .A(_1317_), .B(_1598_), .C(_1600_), .Y(_1229_) );
NAND2X1 NAND2X1_247 ( .A(reg_file_inst_mem_5__2_), .B(_1598_), .Y(_1601_) );
OAI21X1 OAI21X1_322 ( .A(_1319_), .B(_1598_), .C(_1601_), .Y(_1230_) );
NAND2X1 NAND2X1_248 ( .A(reg_file_inst_mem_5__3_), .B(_1598_), .Y(_1602_) );
OAI21X1 OAI21X1_323 ( .A(_1321_), .B(_1598_), .C(_1602_), .Y(_1231_) );
NAND2X1 NAND2X1_249 ( .A(reg_file_inst_mem_5__4_), .B(_1598_), .Y(_1603_) );
OAI21X1 OAI21X1_324 ( .A(_1323_), .B(_1598_), .C(_1603_), .Y(_1232_) );
NAND2X1 NAND2X1_250 ( .A(reg_file_inst_mem_5__5_), .B(_1598_), .Y(_1604_) );
OAI21X1 OAI21X1_325 ( .A(_1325_), .B(_1598_), .C(_1604_), .Y(_1233_) );
NAND2X1 NAND2X1_251 ( .A(reg_file_inst_mem_5__6_), .B(_1598_), .Y(_1605_) );
OAI21X1 OAI21X1_326 ( .A(_1327_), .B(_1598_), .C(_1605_), .Y(_1234_) );
NAND2X1 NAND2X1_252 ( .A(reg_file_inst_mem_5__7_), .B(_1598_), .Y(_1606_) );
OAI21X1 OAI21X1_327 ( .A(_1329_), .B(_1598_), .C(_1606_), .Y(_1235_) );
NAND2X1 NAND2X1_253 ( .A(_1311_), .B(_1371_), .Y(_1607_) );
NAND2X1 NAND2X1_254 ( .A(reg_file_inst_mem_6__0_), .B(_1607_), .Y(_1608_) );
OAI21X1 OAI21X1_328 ( .A(_1308_), .B(_1607_), .C(_1608_), .Y(_1236_) );
NAND2X1 NAND2X1_255 ( .A(reg_file_inst_mem_6__1_), .B(_1607_), .Y(_1609_) );
OAI21X1 OAI21X1_329 ( .A(_1317_), .B(_1607_), .C(_1609_), .Y(_1237_) );
NAND2X1 NAND2X1_256 ( .A(reg_file_inst_mem_6__2_), .B(_1607_), .Y(_1610_) );
OAI21X1 OAI21X1_330 ( .A(_1319_), .B(_1607_), .C(_1610_), .Y(_1238_) );
NAND2X1 NAND2X1_257 ( .A(reg_file_inst_mem_6__3_), .B(_1607_), .Y(_1611_) );
OAI21X1 OAI21X1_331 ( .A(_1321_), .B(_1607_), .C(_1611_), .Y(_1239_) );
NAND2X1 NAND2X1_258 ( .A(reg_file_inst_mem_6__4_), .B(_1607_), .Y(_1612_) );
OAI21X1 OAI21X1_332 ( .A(_1323_), .B(_1607_), .C(_1612_), .Y(_1240_) );
NAND2X1 NAND2X1_259 ( .A(reg_file_inst_mem_6__5_), .B(_1607_), .Y(_1613_) );
OAI21X1 OAI21X1_333 ( .A(_1325_), .B(_1607_), .C(_1613_), .Y(_1241_) );
NAND2X1 NAND2X1_260 ( .A(reg_file_inst_mem_6__6_), .B(_1607_), .Y(_1614_) );
OAI21X1 OAI21X1_334 ( .A(_1327_), .B(_1607_), .C(_1614_), .Y(_1242_) );
NAND2X1 NAND2X1_261 ( .A(reg_file_inst_mem_6__7_), .B(_1607_), .Y(_1615_) );
OAI21X1 OAI21X1_335 ( .A(_1329_), .B(_1607_), .C(_1615_), .Y(_1243_) );
NOR2X1 NOR2X1_214 ( .A(_1310_), .B(_1347_), .Y(_1616_) );
NAND2X1 NAND2X1_262 ( .A(reg_file_inst_wr_data_in_0_), .B(_1616_), .Y(_1617_) );
OAI21X1 OAI21X1_336 ( .A(_1342_), .B(_1616_), .C(_1617_), .Y(_1244_) );
NAND2X1 NAND2X1_263 ( .A(reg_file_inst_wr_data_in_1_), .B(_1616_), .Y(_1618_) );
OAI21X1 OAI21X1_337 ( .A(_1389_), .B(_1616_), .C(_1618_), .Y(_1245_) );
NOR2X1 NOR2X1_215 ( .A(reg_file_inst_mem_7__2_), .B(_1616_), .Y(_1619_) );
AOI21X1 AOI21X1_116 ( .A(_1319_), .B(_1616_), .C(_1619_), .Y(_1246_) );
NOR2X1 NOR2X1_216 ( .A(reg_file_inst_mem_7__3_), .B(_1616_), .Y(_1620_) );
AOI21X1 AOI21X1_117 ( .A(_1321_), .B(_1616_), .C(_1620_), .Y(_1247_) );
NAND2X1 NAND2X1_264 ( .A(reg_file_inst_wr_data_in_4_), .B(_1616_), .Y(_1621_) );
OAI21X1 OAI21X1_338 ( .A(_1464_), .B(_1616_), .C(_1621_), .Y(_1248_) );
NOR2X1 NOR2X1_217 ( .A(reg_file_inst_mem_7__5_), .B(_1616_), .Y(_1622_) );
AOI21X1 AOI21X1_118 ( .A(_1325_), .B(_1616_), .C(_1622_), .Y(_1249_) );
NOR2X1 NOR2X1_218 ( .A(reg_file_inst_mem_7__6_), .B(_1616_), .Y(_1623_) );
AOI21X1 AOI21X1_119 ( .A(_1327_), .B(_1616_), .C(_1623_), .Y(_1250_) );
NAND2X1 NAND2X1_265 ( .A(reg_file_inst_wr_data_in_7_), .B(_1616_), .Y(_1624_) );
OAI21X1 OAI21X1_339 ( .A(_1533_), .B(_1616_), .C(_1624_), .Y(_1251_) );
NAND2X1 NAND2X1_266 ( .A(_1311_), .B(_1430_), .Y(_1625_) );
NAND2X1 NAND2X1_267 ( .A(reg_file_inst_mem_8__0_), .B(_1625_), .Y(_1626_) );
OAI21X1 OAI21X1_340 ( .A(_1308_), .B(_1625_), .C(_1626_), .Y(_1252_) );
NAND2X1 NAND2X1_268 ( .A(reg_file_inst_mem_8__1_), .B(_1625_), .Y(_1627_) );
OAI21X1 OAI21X1_341 ( .A(_1317_), .B(_1625_), .C(_1627_), .Y(_1253_) );
NAND2X1 NAND2X1_269 ( .A(reg_file_inst_mem_8__2_), .B(_1625_), .Y(_1628_) );
OAI21X1 OAI21X1_342 ( .A(_1319_), .B(_1625_), .C(_1628_), .Y(_1254_) );
NAND2X1 NAND2X1_270 ( .A(reg_file_inst_mem_8__3_), .B(_1625_), .Y(_1629_) );
OAI21X1 OAI21X1_343 ( .A(_1321_), .B(_1625_), .C(_1629_), .Y(_1255_) );
NAND2X1 NAND2X1_271 ( .A(reg_file_inst_mem_8__4_), .B(_1625_), .Y(_1630_) );
OAI21X1 OAI21X1_344 ( .A(_1323_), .B(_1625_), .C(_1630_), .Y(_1256_) );
NAND2X1 NAND2X1_272 ( .A(reg_file_inst_mem_8__5_), .B(_1625_), .Y(_1631_) );
OAI21X1 OAI21X1_345 ( .A(_1325_), .B(_1625_), .C(_1631_), .Y(_1257_) );
NAND2X1 NAND2X1_273 ( .A(reg_file_inst_mem_8__6_), .B(_1625_), .Y(_1632_) );
OAI21X1 OAI21X1_346 ( .A(_1327_), .B(_1625_), .C(_1632_), .Y(_1258_) );
NAND2X1 NAND2X1_274 ( .A(reg_file_inst_mem_8__7_), .B(_1625_), .Y(_1633_) );
OAI21X1 OAI21X1_347 ( .A(_1329_), .B(_1625_), .C(_1633_), .Y(_1259_) );
NAND2X1 NAND2X1_275 ( .A(_1311_), .B(_1374_), .Y(_1634_) );
OAI21X1 OAI21X1_348 ( .A(_1310_), .B(_1417_), .C(reg_file_inst_mem_9__0_), .Y(_1635_) );
OAI21X1 OAI21X1_349 ( .A(_1308_), .B(_1634_), .C(_1635_), .Y(_1260_) );
OAI21X1 OAI21X1_350 ( .A(_1310_), .B(_1417_), .C(reg_file_inst_mem_9__1_), .Y(_1636_) );
OAI21X1 OAI21X1_351 ( .A(_1317_), .B(_1634_), .C(_1636_), .Y(_1261_) );
OAI21X1 OAI21X1_352 ( .A(_1310_), .B(_1417_), .C(reg_file_inst_mem_9__2_), .Y(_1637_) );
OAI21X1 OAI21X1_353 ( .A(_1319_), .B(_1634_), .C(_1637_), .Y(_1262_) );
OAI21X1 OAI21X1_354 ( .A(_1310_), .B(_1417_), .C(reg_file_inst_mem_9__3_), .Y(_1638_) );
OAI21X1 OAI21X1_355 ( .A(_1321_), .B(_1634_), .C(_1638_), .Y(_1263_) );
OAI21X1 OAI21X1_356 ( .A(_1310_), .B(_1417_), .C(reg_file_inst_mem_9__4_), .Y(_1639_) );
OAI21X1 OAI21X1_357 ( .A(_1323_), .B(_1634_), .C(_1639_), .Y(_1264_) );
OAI21X1 OAI21X1_358 ( .A(_1310_), .B(_1417_), .C(reg_file_inst_mem_9__5_), .Y(_1640_) );
OAI21X1 OAI21X1_359 ( .A(_1325_), .B(_1634_), .C(_1640_), .Y(_1265_) );
OAI21X1 OAI21X1_360 ( .A(_1310_), .B(_1417_), .C(reg_file_inst_mem_9__6_), .Y(_1641_) );
OAI21X1 OAI21X1_361 ( .A(_1327_), .B(_1634_), .C(_1641_), .Y(_1266_) );
OAI21X1 OAI21X1_362 ( .A(_1310_), .B(_1417_), .C(reg_file_inst_mem_9__7_), .Y(_1642_) );
OAI21X1 OAI21X1_363 ( .A(_1329_), .B(_1634_), .C(_1642_), .Y(_1267_) );
NAND2X1 NAND2X1_276 ( .A(_1311_), .B(_1354_), .Y(_1643_) );
NAND2X1 NAND2X1_277 ( .A(reg_file_inst_mem_10__0_), .B(_1643_), .Y(_1644_) );
OAI21X1 OAI21X1_364 ( .A(_1308_), .B(_1643_), .C(_1644_), .Y(_1268_) );
NAND2X1 NAND2X1_278 ( .A(reg_file_inst_mem_10__1_), .B(_1643_), .Y(_1645_) );
OAI21X1 OAI21X1_365 ( .A(_1317_), .B(_1643_), .C(_1645_), .Y(_1269_) );
NAND2X1 NAND2X1_279 ( .A(reg_file_inst_mem_10__2_), .B(_1643_), .Y(_1646_) );
OAI21X1 OAI21X1_366 ( .A(_1319_), .B(_1643_), .C(_1646_), .Y(_1270_) );
NAND2X1 NAND2X1_280 ( .A(reg_file_inst_mem_10__3_), .B(_1643_), .Y(_1647_) );
OAI21X1 OAI21X1_367 ( .A(_1321_), .B(_1643_), .C(_1647_), .Y(_1271_) );
NAND2X1 NAND2X1_281 ( .A(reg_file_inst_mem_10__4_), .B(_1643_), .Y(_1648_) );
OAI21X1 OAI21X1_368 ( .A(_1323_), .B(_1643_), .C(_1648_), .Y(_1272_) );
NAND2X1 NAND2X1_282 ( .A(reg_file_inst_mem_10__5_), .B(_1643_), .Y(_1649_) );
OAI21X1 OAI21X1_369 ( .A(_1325_), .B(_1643_), .C(_1649_), .Y(_1273_) );
NAND2X1 NAND2X1_283 ( .A(reg_file_inst_mem_10__6_), .B(_1643_), .Y(_1650_) );
OAI21X1 OAI21X1_370 ( .A(_1327_), .B(_1643_), .C(_1650_), .Y(_1274_) );
NAND2X1 NAND2X1_284 ( .A(reg_file_inst_mem_10__7_), .B(_1643_), .Y(_1651_) );
OAI21X1 OAI21X1_371 ( .A(_1329_), .B(_1643_), .C(_1651_), .Y(_1275_) );
AND2X2 AND2X2_46 ( .A(_1362_), .B(_1311_), .Y(_1652_) );
NOR2X1 NOR2X1_219 ( .A(reg_file_inst_mem_11__0_), .B(_1652_), .Y(_1653_) );
AOI21X1 AOI21X1_120 ( .A(_1308_), .B(_1652_), .C(_1653_), .Y(_1276_) );
NOR2X1 NOR2X1_220 ( .A(reg_file_inst_mem_11__1_), .B(_1652_), .Y(_1654_) );
AOI21X1 AOI21X1_121 ( .A(_1317_), .B(_1652_), .C(_1654_), .Y(_1277_) );
NOR2X1 NOR2X1_221 ( .A(reg_file_inst_mem_11__2_), .B(_1652_), .Y(_1655_) );
AOI21X1 AOI21X1_122 ( .A(_1319_), .B(_1652_), .C(_1655_), .Y(_1278_) );
NOR2X1 NOR2X1_222 ( .A(reg_file_inst_mem_11__3_), .B(_1652_), .Y(_1656_) );
AOI21X1 AOI21X1_123 ( .A(_1321_), .B(_1652_), .C(_1656_), .Y(_1279_) );
NOR2X1 NOR2X1_223 ( .A(reg_file_inst_mem_11__4_), .B(_1652_), .Y(_1657_) );
AOI21X1 AOI21X1_124 ( .A(_1323_), .B(_1652_), .C(_1657_), .Y(_1280_) );
NOR2X1 NOR2X1_224 ( .A(reg_file_inst_mem_11__5_), .B(_1652_), .Y(_1658_) );
AOI21X1 AOI21X1_125 ( .A(_1325_), .B(_1652_), .C(_1658_), .Y(_1281_) );
NOR2X1 NOR2X1_225 ( .A(reg_file_inst_mem_11__6_), .B(_1652_), .Y(_1659_) );
AOI21X1 AOI21X1_126 ( .A(_1327_), .B(_1652_), .C(_1659_), .Y(_1282_) );
NOR2X1 NOR2X1_226 ( .A(reg_file_inst_mem_11__7_), .B(_1652_), .Y(_1660_) );
AOI21X1 AOI21X1_127 ( .A(_1329_), .B(_1652_), .C(_1660_), .Y(_1283_) );
NAND2X1 NAND2X1_285 ( .A(_1311_), .B(_1358_), .Y(_1661_) );
OAI21X1 OAI21X1_372 ( .A(_1310_), .B(_1359_), .C(reg_file_inst_mem_12__0_), .Y(_1662_) );
OAI21X1 OAI21X1_373 ( .A(_1308_), .B(_1661_), .C(_1662_), .Y(_1284_) );
OAI21X1 OAI21X1_374 ( .A(_1310_), .B(_1359_), .C(reg_file_inst_mem_12__1_), .Y(_1663_) );
OAI21X1 OAI21X1_375 ( .A(_1317_), .B(_1661_), .C(_1663_), .Y(_1285_) );
OAI21X1 OAI21X1_376 ( .A(_1310_), .B(_1359_), .C(reg_file_inst_mem_12__2_), .Y(_1664_) );
OAI21X1 OAI21X1_377 ( .A(_1319_), .B(_1661_), .C(_1664_), .Y(_1286_) );
OAI21X1 OAI21X1_378 ( .A(_1310_), .B(_1359_), .C(reg_file_inst_mem_12__3_), .Y(_1665_) );
OAI21X1 OAI21X1_379 ( .A(_1321_), .B(_1661_), .C(_1665_), .Y(_1287_) );
OAI21X1 OAI21X1_380 ( .A(_1310_), .B(_1359_), .C(reg_file_inst_mem_12__4_), .Y(_1666_) );
OAI21X1 OAI21X1_381 ( .A(_1323_), .B(_1661_), .C(_1666_), .Y(_1288_) );
OAI21X1 OAI21X1_382 ( .A(_1310_), .B(_1359_), .C(reg_file_inst_mem_12__5_), .Y(_1667_) );
OAI21X1 OAI21X1_383 ( .A(_1325_), .B(_1661_), .C(_1667_), .Y(_1289_) );
OAI21X1 OAI21X1_384 ( .A(_1310_), .B(_1359_), .C(reg_file_inst_mem_12__6_), .Y(_1668_) );
OAI21X1 OAI21X1_385 ( .A(_1327_), .B(_1661_), .C(_1668_), .Y(_1290_) );
OAI21X1 OAI21X1_386 ( .A(_1310_), .B(_1359_), .C(reg_file_inst_mem_12__7_), .Y(_1669_) );
OAI21X1 OAI21X1_387 ( .A(_1329_), .B(_1661_), .C(_1669_), .Y(_1291_) );
NOR2X1 NOR2X1_227 ( .A(_1310_), .B(_1349_), .Y(_1670_) );
NAND2X1 NAND2X1_286 ( .A(reg_file_inst_wr_data_in_0_), .B(_1670_), .Y(_1671_) );
OAI21X1 OAI21X1_388 ( .A(_1341_), .B(_1670_), .C(_1671_), .Y(_1292_) );
NAND2X1 NAND2X1_287 ( .A(reg_file_inst_wr_data_in_1_), .B(_1670_), .Y(_1672_) );
OAI21X1 OAI21X1_389 ( .A(_1388_), .B(_1670_), .C(_1672_), .Y(_1293_) );
NOR2X1 NOR2X1_228 ( .A(reg_file_inst_mem_13__2_), .B(_1670_), .Y(_1673_) );
AOI21X1 AOI21X1_128 ( .A(_1319_), .B(_1670_), .C(_1673_), .Y(_1294_) );
NOR2X1 NOR2X1_229 ( .A(reg_file_inst_mem_13__3_), .B(_1670_), .Y(_1674_) );
AOI21X1 AOI21X1_129 ( .A(_1321_), .B(_1670_), .C(_1674_), .Y(_1295_) );
NAND2X1 NAND2X1_288 ( .A(reg_file_inst_wr_data_in_4_), .B(_1670_), .Y(_1675_) );
OAI21X1 OAI21X1_390 ( .A(_1463_), .B(_1670_), .C(_1675_), .Y(_1296_) );
NOR2X1 NOR2X1_230 ( .A(reg_file_inst_mem_13__5_), .B(_1670_), .Y(_1676_) );
AOI21X1 AOI21X1_130 ( .A(_1325_), .B(_1670_), .C(_1676_), .Y(_1297_) );
NOR2X1 NOR2X1_231 ( .A(reg_file_inst_mem_13__6_), .B(_1670_), .Y(_1677_) );
AOI21X1 AOI21X1_131 ( .A(_1327_), .B(_1670_), .C(_1677_), .Y(_1298_) );
NAND2X1 NAND2X1_289 ( .A(reg_file_inst_wr_data_in_7_), .B(_1670_), .Y(_1678_) );
OAI21X1 OAI21X1_391 ( .A(_1532_), .B(_1670_), .C(_1678_), .Y(_1299_) );
NOR2X1 NOR2X1_232 ( .A(_1310_), .B(_1410_), .Y(_1679_) );
NOR2X1 NOR2X1_233 ( .A(reg_file_inst_mem_14__0_), .B(_1679_), .Y(_1680_) );
AOI21X1 AOI21X1_132 ( .A(_1308_), .B(_1679_), .C(_1680_), .Y(_1300_) );
NOR2X1 NOR2X1_234 ( .A(reg_file_inst_mem_14__1_), .B(_1679_), .Y(_1681_) );
AOI21X1 AOI21X1_133 ( .A(_1317_), .B(_1679_), .C(_1681_), .Y(_1301_) );
NAND2X1 NAND2X1_290 ( .A(reg_file_inst_wr_data_in_2_), .B(_1679_), .Y(_1682_) );
OAI21X1 OAI21X1_392 ( .A(_1409_), .B(_1679_), .C(_1682_), .Y(_1302_) );
NAND2X1 NAND2X1_291 ( .A(reg_file_inst_wr_data_in_3_), .B(_1679_), .Y(_1683_) );
OAI21X1 OAI21X1_393 ( .A(_1438_), .B(_1679_), .C(_1683_), .Y(_1303_) );
NOR2X1 NOR2X1_235 ( .A(reg_file_inst_mem_14__4_), .B(_1679_), .Y(_1684_) );
AOI21X1 AOI21X1_134 ( .A(_1323_), .B(_1679_), .C(_1684_), .Y(_1304_) );
NAND2X1 NAND2X1_292 ( .A(reg_file_inst_wr_data_in_5_), .B(_1679_), .Y(_1685_) );
OAI21X1 OAI21X1_394 ( .A(_1484_), .B(_1679_), .C(_1685_), .Y(_1305_) );
NAND2X1 NAND2X1_293 ( .A(reg_file_inst_wr_data_in_6_), .B(_1679_), .Y(_1686_) );
OAI21X1 OAI21X1_395 ( .A(_1507_), .B(_1679_), .C(_1686_), .Y(_1306_) );
NOR2X1 NOR2X1_236 ( .A(reg_file_inst_mem_14__7_), .B(_1679_), .Y(_1687_) );
AOI21X1 AOI21X1_135 ( .A(_1329_), .B(_1679_), .C(_1687_), .Y(_1307_) );
INVX1 INVX1_243 ( .A(reg_file_inst_rd_data_valid_out), .Y(_1688_) );
OAI21X1 OAI21X1_396 ( .A(_1688_), .B(_1310_), .C(_1333_), .Y(_1187_) );
DFFSR DFFSR_50 ( .CLK(ref_clk), .D(_1171_), .Q(reg_file_inst_mem_15__0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_51 ( .CLK(ref_clk), .D(_1172_), .Q(reg_file_inst_mem_15__1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_52 ( .CLK(ref_clk), .D(_1173_), .Q(reg_file_inst_mem_15__2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_53 ( .CLK(ref_clk), .D(_1174_), .Q(reg_file_inst_mem_15__3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_54 ( .CLK(ref_clk), .D(_1175_), .Q(reg_file_inst_mem_15__4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_55 ( .CLK(ref_clk), .D(_1176_), .Q(reg_file_inst_mem_15__5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_56 ( .CLK(ref_clk), .D(_1177_), .Q(reg_file_inst_mem_15__6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_57 ( .CLK(ref_clk), .D(_1178_), .Q(reg_file_inst_mem_15__7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_58 ( .CLK(ref_clk), .D(_1179_), .Q(reg_file_inst_rd_data_out_0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_59 ( .CLK(ref_clk), .D(_1180_), .Q(reg_file_inst_rd_data_out_1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_60 ( .CLK(ref_clk), .D(_1181_), .Q(reg_file_inst_rd_data_out_2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_61 ( .CLK(ref_clk), .D(_1182_), .Q(reg_file_inst_rd_data_out_3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_62 ( .CLK(ref_clk), .D(_1183_), .Q(reg_file_inst_rd_data_out_4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_63 ( .CLK(ref_clk), .D(_1184_), .Q(reg_file_inst_rd_data_out_5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_64 ( .CLK(ref_clk), .D(_1185_), .Q(reg_file_inst_rd_data_out_6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_65 ( .CLK(ref_clk), .D(_1186_), .Q(reg_file_inst_rd_data_out_7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_66 ( .CLK(ref_clk), .D(_1187_), .Q(reg_file_inst_rd_data_valid_out), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_67 ( .CLK(ref_clk), .D(_1188_), .Q(alu_inst_data_a_in_0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_68 ( .CLK(ref_clk), .D(_1189_), .Q(alu_inst_data_a_in_1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_69 ( .CLK(ref_clk), .D(_1190_), .Q(alu_inst_data_a_in_2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_70 ( .CLK(ref_clk), .D(_1191_), .Q(alu_inst_data_a_in_3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_71 ( .CLK(ref_clk), .D(_1192_), .Q(alu_inst_data_a_in_4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_72 ( .CLK(ref_clk), .D(_1193_), .Q(alu_inst_data_a_in_5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_73 ( .CLK(ref_clk), .D(_1194_), .Q(alu_inst_data_a_in_6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_74 ( .CLK(ref_clk), .D(_1195_), .Q(alu_inst_data_a_in_7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_75 ( .CLK(ref_clk), .D(_1196_), .Q(alu_inst_data_b_in_0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_76 ( .CLK(ref_clk), .D(_1197_), .Q(alu_inst_data_b_in_1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_77 ( .CLK(ref_clk), .D(_1198_), .Q(alu_inst_data_b_in_2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_78 ( .CLK(ref_clk), .D(_1199_), .Q(alu_inst_data_b_in_3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_79 ( .CLK(ref_clk), .D(_1200_), .Q(alu_inst_data_b_in_4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_80 ( .CLK(ref_clk), .D(_1201_), .Q(alu_inst_data_b_in_5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_81 ( .CLK(ref_clk), .D(_1202_), .Q(alu_inst_data_b_in_6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_82 ( .CLK(ref_clk), .D(_1203_), .Q(alu_inst_data_b_in_7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_83 ( .CLK(ref_clk), .D(_1204_), .Q(uart_top_inst_par_en_in), .R(_true), .S(alu_inst_reset_n) );
DFFSR DFFSR_84 ( .CLK(ref_clk), .D(_1205_), .Q(uart_top_inst_par_type_in), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_85 ( .CLK(ref_clk), .D(_1206_), .Q(reg_file_inst_mem_2__2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_86 ( .CLK(ref_clk), .D(_1207_), .Q(reg_file_inst_mem_2__3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_87 ( .CLK(ref_clk), .D(_1208_), .Q(reg_file_inst_mem_2__4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_88 ( .CLK(ref_clk), .D(_1209_), .Q(reg_file_inst_mem_2__5_), .R(_true), .S(alu_inst_reset_n) );
DFFSR DFFSR_89 ( .CLK(ref_clk), .D(_1210_), .Q(reg_file_inst_mem_2__6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_90 ( .CLK(ref_clk), .D(_1211_), .Q(reg_file_inst_mem_2__7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_91 ( .CLK(ref_clk), .D(_1212_), .Q(clk_divider_inst_div_ratio_in_0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_92 ( .CLK(ref_clk), .D(_1213_), .Q(clk_divider_inst_div_ratio_in_1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_93 ( .CLK(ref_clk), .D(_1214_), .Q(clk_divider_inst_div_ratio_in_2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_94 ( .CLK(ref_clk), .D(_1215_), .Q(clk_divider_inst_div_ratio_in_3_), .R(_true), .S(alu_inst_reset_n) );
DFFSR DFFSR_95 ( .CLK(ref_clk), .D(_1216_), .Q(clk_divider_inst_div_ratio_in_4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_96 ( .CLK(ref_clk), .D(_1217_), .Q(reg_file_inst_mem_3__5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_97 ( .CLK(ref_clk), .D(_1218_), .Q(reg_file_inst_mem_3__6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_98 ( .CLK(ref_clk), .D(_1219_), .Q(reg_file_inst_mem_3__7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_99 ( .CLK(ref_clk), .D(_1220_), .Q(reg_file_inst_mem_4__0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_100 ( .CLK(ref_clk), .D(_1221_), .Q(reg_file_inst_mem_4__1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_101 ( .CLK(ref_clk), .D(_1222_), .Q(reg_file_inst_mem_4__2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_102 ( .CLK(ref_clk), .D(_1223_), .Q(reg_file_inst_mem_4__3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_103 ( .CLK(ref_clk), .D(_1224_), .Q(reg_file_inst_mem_4__4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_104 ( .CLK(ref_clk), .D(_1225_), .Q(reg_file_inst_mem_4__5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_105 ( .CLK(ref_clk), .D(_1226_), .Q(reg_file_inst_mem_4__6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_106 ( .CLK(ref_clk), .D(_1227_), .Q(reg_file_inst_mem_4__7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_107 ( .CLK(ref_clk), .D(_1228_), .Q(reg_file_inst_mem_5__0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_108 ( .CLK(ref_clk), .D(_1229_), .Q(reg_file_inst_mem_5__1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_109 ( .CLK(ref_clk), .D(_1230_), .Q(reg_file_inst_mem_5__2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_110 ( .CLK(ref_clk), .D(_1231_), .Q(reg_file_inst_mem_5__3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_111 ( .CLK(ref_clk), .D(_1232_), .Q(reg_file_inst_mem_5__4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_112 ( .CLK(ref_clk), .D(_1233_), .Q(reg_file_inst_mem_5__5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_113 ( .CLK(ref_clk), .D(_1234_), .Q(reg_file_inst_mem_5__6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_114 ( .CLK(ref_clk), .D(_1235_), .Q(reg_file_inst_mem_5__7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_115 ( .CLK(ref_clk), .D(_1236_), .Q(reg_file_inst_mem_6__0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_116 ( .CLK(ref_clk), .D(_1237_), .Q(reg_file_inst_mem_6__1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_117 ( .CLK(ref_clk), .D(_1238_), .Q(reg_file_inst_mem_6__2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_118 ( .CLK(ref_clk), .D(_1239_), .Q(reg_file_inst_mem_6__3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_119 ( .CLK(ref_clk), .D(_1240_), .Q(reg_file_inst_mem_6__4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_120 ( .CLK(ref_clk), .D(_1241_), .Q(reg_file_inst_mem_6__5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_121 ( .CLK(ref_clk), .D(_1242_), .Q(reg_file_inst_mem_6__6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_122 ( .CLK(ref_clk), .D(_1243_), .Q(reg_file_inst_mem_6__7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_123 ( .CLK(ref_clk), .D(_1244_), .Q(reg_file_inst_mem_7__0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_124 ( .CLK(ref_clk), .D(_1245_), .Q(reg_file_inst_mem_7__1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_125 ( .CLK(ref_clk), .D(_1246_), .Q(reg_file_inst_mem_7__2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_126 ( .CLK(ref_clk), .D(_1247_), .Q(reg_file_inst_mem_7__3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_127 ( .CLK(ref_clk), .D(_1248_), .Q(reg_file_inst_mem_7__4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_128 ( .CLK(ref_clk), .D(_1249_), .Q(reg_file_inst_mem_7__5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_129 ( .CLK(ref_clk), .D(_1250_), .Q(reg_file_inst_mem_7__6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_130 ( .CLK(ref_clk), .D(_1251_), .Q(reg_file_inst_mem_7__7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_131 ( .CLK(ref_clk), .D(_1252_), .Q(reg_file_inst_mem_8__0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_132 ( .CLK(ref_clk), .D(_1253_), .Q(reg_file_inst_mem_8__1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_133 ( .CLK(ref_clk), .D(_1254_), .Q(reg_file_inst_mem_8__2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_134 ( .CLK(ref_clk), .D(_1255_), .Q(reg_file_inst_mem_8__3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_135 ( .CLK(ref_clk), .D(_1256_), .Q(reg_file_inst_mem_8__4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_136 ( .CLK(ref_clk), .D(_1257_), .Q(reg_file_inst_mem_8__5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_137 ( .CLK(ref_clk), .D(_1258_), .Q(reg_file_inst_mem_8__6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_138 ( .CLK(ref_clk), .D(_1259_), .Q(reg_file_inst_mem_8__7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_139 ( .CLK(ref_clk), .D(_1260_), .Q(reg_file_inst_mem_9__0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_140 ( .CLK(ref_clk), .D(_1261_), .Q(reg_file_inst_mem_9__1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_141 ( .CLK(ref_clk), .D(_1262_), .Q(reg_file_inst_mem_9__2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_142 ( .CLK(ref_clk), .D(_1263_), .Q(reg_file_inst_mem_9__3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_143 ( .CLK(ref_clk), .D(_1264_), .Q(reg_file_inst_mem_9__4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_144 ( .CLK(ref_clk), .D(_1265_), .Q(reg_file_inst_mem_9__5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_145 ( .CLK(ref_clk), .D(_1266_), .Q(reg_file_inst_mem_9__6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_146 ( .CLK(ref_clk), .D(_1267_), .Q(reg_file_inst_mem_9__7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_147 ( .CLK(ref_clk), .D(_1268_), .Q(reg_file_inst_mem_10__0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_148 ( .CLK(ref_clk), .D(_1269_), .Q(reg_file_inst_mem_10__1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_149 ( .CLK(ref_clk), .D(_1270_), .Q(reg_file_inst_mem_10__2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_150 ( .CLK(ref_clk), .D(_1271_), .Q(reg_file_inst_mem_10__3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_151 ( .CLK(ref_clk), .D(_1272_), .Q(reg_file_inst_mem_10__4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_152 ( .CLK(ref_clk), .D(_1273_), .Q(reg_file_inst_mem_10__5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_153 ( .CLK(ref_clk), .D(_1274_), .Q(reg_file_inst_mem_10__6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_154 ( .CLK(ref_clk), .D(_1275_), .Q(reg_file_inst_mem_10__7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_155 ( .CLK(ref_clk), .D(_1276_), .Q(reg_file_inst_mem_11__0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_156 ( .CLK(ref_clk), .D(_1277_), .Q(reg_file_inst_mem_11__1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_157 ( .CLK(ref_clk), .D(_1278_), .Q(reg_file_inst_mem_11__2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_158 ( .CLK(ref_clk), .D(_1279_), .Q(reg_file_inst_mem_11__3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_159 ( .CLK(ref_clk), .D(_1280_), .Q(reg_file_inst_mem_11__4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_160 ( .CLK(ref_clk), .D(_1281_), .Q(reg_file_inst_mem_11__5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_161 ( .CLK(ref_clk), .D(_1282_), .Q(reg_file_inst_mem_11__6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_162 ( .CLK(ref_clk), .D(_1283_), .Q(reg_file_inst_mem_11__7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_163 ( .CLK(ref_clk), .D(_1284_), .Q(reg_file_inst_mem_12__0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_164 ( .CLK(ref_clk), .D(_1285_), .Q(reg_file_inst_mem_12__1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_165 ( .CLK(ref_clk), .D(_1286_), .Q(reg_file_inst_mem_12__2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_166 ( .CLK(ref_clk), .D(_1287_), .Q(reg_file_inst_mem_12__3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_167 ( .CLK(ref_clk), .D(_1288_), .Q(reg_file_inst_mem_12__4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_168 ( .CLK(ref_clk), .D(_1289_), .Q(reg_file_inst_mem_12__5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_169 ( .CLK(ref_clk), .D(_1290_), .Q(reg_file_inst_mem_12__6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_170 ( .CLK(ref_clk), .D(_1291_), .Q(reg_file_inst_mem_12__7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_171 ( .CLK(ref_clk), .D(_1292_), .Q(reg_file_inst_mem_13__0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_172 ( .CLK(ref_clk), .D(_1293_), .Q(reg_file_inst_mem_13__1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_173 ( .CLK(ref_clk), .D(_1294_), .Q(reg_file_inst_mem_13__2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_174 ( .CLK(ref_clk), .D(_1295_), .Q(reg_file_inst_mem_13__3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_175 ( .CLK(ref_clk), .D(_1296_), .Q(reg_file_inst_mem_13__4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_176 ( .CLK(ref_clk), .D(_1297_), .Q(reg_file_inst_mem_13__5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_177 ( .CLK(ref_clk), .D(_1298_), .Q(reg_file_inst_mem_13__6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_178 ( .CLK(ref_clk), .D(_1299_), .Q(reg_file_inst_mem_13__7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_179 ( .CLK(ref_clk), .D(_1300_), .Q(reg_file_inst_mem_14__0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_180 ( .CLK(ref_clk), .D(_1301_), .Q(reg_file_inst_mem_14__1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_181 ( .CLK(ref_clk), .D(_1302_), .Q(reg_file_inst_mem_14__2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_182 ( .CLK(ref_clk), .D(_1303_), .Q(reg_file_inst_mem_14__3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_183 ( .CLK(ref_clk), .D(_1304_), .Q(reg_file_inst_mem_14__4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_184 ( .CLK(ref_clk), .D(_1305_), .Q(reg_file_inst_mem_14__5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_185 ( .CLK(ref_clk), .D(_1306_), .Q(reg_file_inst_mem_14__6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_186 ( .CLK(ref_clk), .D(_1307_), .Q(reg_file_inst_mem_14__7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_187 ( .CLK(ref_clk), .D(reset_synchronizer_inst_0_ff_1_), .Q(alu_inst_reset_n), .R(reset_n), .S(_true) );
DFFSR DFFSR_188 ( .CLK(ref_clk), .D(reset_synchronizer_inst_0_ff_2_), .Q(reset_synchronizer_inst_0_ff_1_), .R(reset_n), .S(_true) );
DFFSR DFFSR_189 ( .CLK(ref_clk), .D(_true), .Q(reset_synchronizer_inst_0_ff_2_), .R(reset_n), .S(_true) );
DFFSR DFFSR_190 ( .CLK(uart_clk), .D(reset_synchronizer_inst_1_ff_1_), .Q(clk_divider_inst_reset_n), .R(reset_n), .S(_true) );
DFFSR DFFSR_191 ( .CLK(uart_clk), .D(reset_synchronizer_inst_1_ff_2_), .Q(reset_synchronizer_inst_1_ff_1_), .R(reset_n), .S(_true) );
DFFSR DFFSR_192 ( .CLK(uart_clk), .D(_true), .Q(reset_synchronizer_inst_1_ff_2_), .R(reset_n), .S(_true) );
INVX1 INVX1_244 ( .A(sys_control_inst_sys_control_rx_inst_current_state_0_), .Y(_1718_) );
NAND2X1 NAND2X1_294 ( .A(sys_control_inst_sys_control_rx_inst_current_state_1_), .B(_1718_), .Y(_1719_) );
INVX1 INVX1_245 ( .A(sys_control_inst_sys_control_rx_inst_current_state_3_), .Y(_1720_) );
NAND2X1 NAND2X1_295 ( .A(sys_control_inst_sys_control_rx_inst_current_state_2_), .B(_1720_), .Y(_1721_) );
NOR2X1 NOR2X1_237 ( .A(_1719_), .B(_1721_), .Y(reg_file_inst_rd_en_in) );
INVX1 INVX1_246 ( .A(data_synchronizer_inst_0_enable_pulse_out), .Y(_1722_) );
INVX1 INVX1_247 ( .A(sys_control_inst_sys_control_rx_inst_current_state_2_), .Y(_1723_) );
NAND2X1 NAND2X1_296 ( .A(sys_control_inst_sys_control_rx_inst_current_state_3_), .B(_1723_), .Y(_1724_) );
INVX1 INVX1_248 ( .A(sys_control_inst_sys_control_rx_inst_current_state_1_), .Y(_1725_) );
NAND2X1 NAND2X1_297 ( .A(sys_control_inst_sys_control_rx_inst_current_state_0_), .B(_1725_), .Y(_1726_) );
NOR2X1 NOR2X1_238 ( .A(_1724_), .B(_1726_), .Y(_1727_) );
INVX1 INVX1_249 ( .A(_1727_), .Y(_1728_) );
NOR2X1 NOR2X1_239 ( .A(_1722_), .B(_1728_), .Y(alu_inst_alu_out_comp_valid) );
OAI21X1 OAI21X1_397 ( .A(_1719_), .B(_1724_), .C(_1728_), .Y(clk_gate_inst_clk_en_in) );
AND2X2 AND2X2_47 ( .A(_1727_), .B(data_synchronizer_inst_0_sync_data_out_0_), .Y(alu_inst_alu_func_in_0_) );
AND2X2 AND2X2_48 ( .A(_1727_), .B(data_synchronizer_inst_0_sync_data_out_1_), .Y(alu_inst_alu_func_in_1_) );
AND2X2 AND2X2_49 ( .A(_1727_), .B(data_synchronizer_inst_0_sync_data_out_2_), .Y(alu_inst_alu_func_in_2_) );
AND2X2 AND2X2_50 ( .A(_1727_), .B(data_synchronizer_inst_0_sync_data_out_3_), .Y(alu_inst_alu_func_in_3_) );
INVX1 INVX1_250 ( .A(sys_control_inst_sys_control_rx_inst_rf_addr_reg_0_), .Y(_1729_) );
NOR2X1 NOR2X1_240 ( .A(sys_control_inst_sys_control_rx_inst_current_state_3_), .B(sys_control_inst_sys_control_rx_inst_current_state_2_), .Y(_1730_) );
AND2X2 AND2X2_51 ( .A(sys_control_inst_sys_control_rx_inst_current_state_1_), .B(sys_control_inst_sys_control_rx_inst_current_state_0_), .Y(_1731_) );
AOI21X1 AOI21X1_136 ( .A(_1730_), .B(_1731_), .C(reg_file_inst_rd_en_in), .Y(_1732_) );
NOR2X1 NOR2X1_241 ( .A(sys_control_inst_sys_control_rx_inst_current_state_2_), .B(_1720_), .Y(_1733_) );
NOR2X1 NOR2X1_242 ( .A(sys_control_inst_sys_control_rx_inst_current_state_1_), .B(sys_control_inst_sys_control_rx_inst_current_state_0_), .Y(_1734_) );
AND2X2 AND2X2_52 ( .A(_1733_), .B(_1734_), .Y(_1735_) );
INVX1 INVX1_251 ( .A(_1735_), .Y(_1736_) );
OAI21X1 OAI21X1_398 ( .A(_1729_), .B(_1732_), .C(_1736_), .Y(reg_file_inst_addr_in_0_) );
INVX1 INVX1_252 ( .A(sys_control_inst_sys_control_rx_inst_rf_addr_reg_1_), .Y(_1737_) );
NOR2X1 NOR2X1_243 ( .A(_1737_), .B(_1732_), .Y(reg_file_inst_addr_in_1_) );
INVX1 INVX1_253 ( .A(sys_control_inst_sys_control_rx_inst_rf_addr_reg_2_), .Y(_1738_) );
NOR2X1 NOR2X1_244 ( .A(_1738_), .B(_1732_), .Y(reg_file_inst_addr_in_2_) );
INVX1 INVX1_254 ( .A(sys_control_inst_sys_control_rx_inst_rf_addr_reg_3_), .Y(_1739_) );
NOR2X1 NOR2X1_245 ( .A(_1739_), .B(_1732_), .Y(reg_file_inst_addr_in_3_) );
NOR2X1 NOR2X1_246 ( .A(data_synchronizer_inst_0_sync_data_out_2_), .B(data_synchronizer_inst_0_sync_data_out_6_), .Y(_1740_) );
NAND3X1 NAND3X1_202 ( .A(data_synchronizer_inst_0_sync_data_out_3_), .B(data_synchronizer_inst_0_sync_data_out_7_), .C(_1740_), .Y(_1741_) );
NAND2X1 NAND2X1_298 ( .A(data_synchronizer_inst_0_sync_data_out_0_), .B(data_synchronizer_inst_0_sync_data_out_4_), .Y(_1742_) );
INVX1 INVX1_255 ( .A(_1742_), .Y(_1743_) );
NAND3X1 NAND3X1_203 ( .A(data_synchronizer_inst_0_sync_data_out_1_), .B(data_synchronizer_inst_0_sync_data_out_5_), .C(_1743_), .Y(_1744_) );
AND2X2 AND2X2_53 ( .A(data_synchronizer_inst_0_sync_data_out_2_), .B(data_synchronizer_inst_0_sync_data_out_3_), .Y(_1745_) );
NOR2X1 NOR2X1_247 ( .A(data_synchronizer_inst_0_sync_data_out_1_), .B(data_synchronizer_inst_0_sync_data_out_5_), .Y(_1746_) );
NAND2X1 NAND2X1_299 ( .A(_1746_), .B(_1745_), .Y(_1747_) );
NOR2X1 NOR2X1_248 ( .A(data_synchronizer_inst_0_sync_data_out_0_), .B(data_synchronizer_inst_0_sync_data_out_4_), .Y(_1748_) );
AND2X2 AND2X2_54 ( .A(data_synchronizer_inst_0_sync_data_out_7_), .B(data_synchronizer_inst_0_sync_data_out_6_), .Y(_1749_) );
NAND2X1 NAND2X1_300 ( .A(_1748_), .B(_1749_), .Y(_1750_) );
OAI22X1 OAI22X1_10 ( .A(_1747_), .B(_1750_), .C(_1741_), .D(_1744_), .Y(_1751_) );
NAND3X1 NAND3X1_204 ( .A(data_synchronizer_inst_0_enable_pulse_out), .B(_1730_), .C(_1734_), .Y(_1752_) );
INVX1 INVX1_256 ( .A(_1752_), .Y(_1753_) );
NAND2X1 NAND2X1_301 ( .A(_1753_), .B(_1751_), .Y(_1754_) );
NOR2X1 NOR2X1_249 ( .A(_1721_), .B(_1726_), .Y(_1755_) );
OAI21X1 OAI21X1_399 ( .A(_1724_), .B(_1726_), .C(_1722_), .Y(_1756_) );
OAI22X1 OAI22X1_11 ( .A(_1755_), .B(_1756_), .C(_1722_), .D(_1735_), .Y(_1757_) );
NAND2X1 NAND2X1_302 ( .A(data_synchronizer_inst_0_enable_pulse_out), .B(_1745_), .Y(_1758_) );
NOR2X1 NOR2X1_250 ( .A(_1742_), .B(_1758_), .Y(_1759_) );
NAND2X1 NAND2X1_303 ( .A(_1746_), .B(_1749_), .Y(_1760_) );
NAND2X1 NAND2X1_304 ( .A(_1730_), .B(_1734_), .Y(_1761_) );
NOR2X1 NOR2X1_251 ( .A(_1760_), .B(_1761_), .Y(_1762_) );
NAND3X1 NAND3X1_205 ( .A(sys_control_inst_sys_control_rx_inst_current_state_1_), .B(_1718_), .C(_1730_), .Y(_1763_) );
NAND2X1 NAND2X1_305 ( .A(_1720_), .B(_1731_), .Y(_1764_) );
MUX2X1 MUX2X1_2 ( .A(_1763_), .B(_1764_), .S(data_synchronizer_inst_0_enable_pulse_out), .Y(_1765_) );
AOI21X1 AOI21X1_137 ( .A(_1762_), .B(_1759_), .C(_1765_), .Y(_1766_) );
NAND3X1 NAND3X1_206 ( .A(_1757_), .B(_1766_), .C(_1754_), .Y(sys_control_inst_sys_control_rx_inst_next_state_0_) );
NOR2X1 NOR2X1_252 ( .A(sys_control_inst_sys_control_rx_inst_current_state_0_), .B(_1725_), .Y(_1767_) );
AOI22X1 AOI22X1_46 ( .A(_1767_), .B(_1730_), .C(_1727_), .D(data_synchronizer_inst_0_enable_pulse_out), .Y(_1768_) );
INVX1 INVX1_257 ( .A(_1764_), .Y(_1769_) );
NAND3X1 NAND3X1_207 ( .A(data_synchronizer_inst_0_sync_data_out_1_), .B(data_synchronizer_inst_0_sync_data_out_5_), .C(_1748_), .Y(_1770_) );
OAI22X1 OAI22X1_12 ( .A(_1747_), .B(_1750_), .C(_1741_), .D(_1770_), .Y(_1771_) );
AOI22X1 AOI22X1_47 ( .A(_1722_), .B(_1769_), .C(_1771_), .D(_1753_), .Y(_1772_) );
NOR2X1 NOR2X1_253 ( .A(sys_control_inst_sys_control_rx_inst_current_state_3_), .B(_1723_), .Y(_1773_) );
NOR2X1 NOR2X1_254 ( .A(sys_control_inst_sys_control_rx_inst_current_state_1_), .B(_1718_), .Y(_1774_) );
NAND3X1 NAND3X1_208 ( .A(data_synchronizer_inst_0_enable_pulse_out), .B(_1773_), .C(_1774_), .Y(_1775_) );
INVX1 INVX1_258 ( .A(reg_file_inst_rd_data_valid_out), .Y(_1776_) );
NAND3X1 NAND3X1_209 ( .A(_1776_), .B(_1767_), .C(_1773_), .Y(_1777_) );
INVX1 INVX1_259 ( .A(alu_inst_data_valid_out), .Y(_1778_) );
NAND3X1 NAND3X1_210 ( .A(_1778_), .B(_1767_), .C(_1733_), .Y(_1779_) );
NAND3X1 NAND3X1_211 ( .A(_1775_), .B(_1777_), .C(_1779_), .Y(_1780_) );
INVX1 INVX1_260 ( .A(_1780_), .Y(_1781_) );
NAND3X1 NAND3X1_212 ( .A(_1768_), .B(_1772_), .C(_1781_), .Y(sys_control_inst_sys_control_rx_inst_next_state_1_) );
NOR2X1 NOR2X1_255 ( .A(_1723_), .B(_1764_), .Y(_1782_) );
AOI21X1 AOI21X1_138 ( .A(_1782_), .B(_1722_), .C(_1755_), .Y(_1783_) );
NAND3X1 NAND3X1_213 ( .A(_1777_), .B(_1783_), .C(_1754_), .Y(sys_control_inst_sys_control_rx_inst_next_state_2_) );
NAND2X1 NAND2X1_306 ( .A(_1759_), .B(_1762_), .Y(_1784_) );
NAND2X1 NAND2X1_307 ( .A(data_synchronizer_inst_0_enable_pulse_out), .B(_1782_), .Y(_1785_) );
NOR2X1 NOR2X1_256 ( .A(_1719_), .B(_1724_), .Y(_1786_) );
AOI22X1 AOI22X1_48 ( .A(_1725_), .B(_1733_), .C(_1786_), .D(_1778_), .Y(_1787_) );
NAND3X1 NAND3X1_214 ( .A(_1787_), .B(_1785_), .C(_1784_), .Y(sys_control_inst_sys_control_rx_inst_next_state_3_) );
NAND2X1 NAND2X1_308 ( .A(alu_inst_data_valid_out), .B(_1786_), .Y(_1788_) );
INVX1 INVX1_261 ( .A(_1788_), .Y(sys_control_inst_sys_control_rx_inst_alu_data_store) );
NAND2X1 NAND2X1_309 ( .A(reg_file_inst_rd_data_valid_out), .B(reg_file_inst_rd_en_in), .Y(_1789_) );
INVX1 INVX1_262 ( .A(_1789_), .Y(sys_control_inst_sys_control_rx_inst_rf_rd_store) );
NOR2X1 NOR2X1_257 ( .A(_1769_), .B(_1735_), .Y(_1689_) );
NOR2X1 NOR2X1_258 ( .A(_1722_), .B(_1689_), .Y(reg_file_inst_wr_en_in) );
OAI21X1 OAI21X1_400 ( .A(_1722_), .B(_1763_), .C(_1775_), .Y(_1790_) );
NAND2X1 NAND2X1_310 ( .A(data_synchronizer_inst_0_sync_data_out_0_), .B(_1790_), .Y(_1791_) );
OAI21X1 OAI21X1_401 ( .A(_1729_), .B(_1790_), .C(_1791_), .Y(_1690_) );
NAND2X1 NAND2X1_311 ( .A(data_synchronizer_inst_0_sync_data_out_1_), .B(_1790_), .Y(_1792_) );
OAI21X1 OAI21X1_402 ( .A(_1737_), .B(_1790_), .C(_1792_), .Y(_1691_) );
NAND2X1 NAND2X1_312 ( .A(data_synchronizer_inst_0_sync_data_out_2_), .B(_1790_), .Y(_1793_) );
OAI21X1 OAI21X1_403 ( .A(_1738_), .B(_1790_), .C(_1793_), .Y(_1692_) );
NAND2X1 NAND2X1_313 ( .A(data_synchronizer_inst_0_sync_data_out_3_), .B(_1790_), .Y(_1794_) );
OAI21X1 OAI21X1_404 ( .A(_1739_), .B(_1790_), .C(_1794_), .Y(_1693_) );
INVX1 INVX1_263 ( .A(alu_inst_data_out_0_), .Y(_1795_) );
NAND2X1 NAND2X1_314 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_0_), .B(_1788_), .Y(_1796_) );
OAI21X1 OAI21X1_405 ( .A(_1795_), .B(_1788_), .C(_1796_), .Y(_1694_) );
INVX1 INVX1_264 ( .A(alu_inst_data_out_1_), .Y(_1797_) );
NAND2X1 NAND2X1_315 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_1_), .B(_1788_), .Y(_1798_) );
OAI21X1 OAI21X1_406 ( .A(_1797_), .B(_1788_), .C(_1798_), .Y(_1695_) );
INVX1 INVX1_265 ( .A(alu_inst_data_out_2_), .Y(_1799_) );
NAND2X1 NAND2X1_316 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_2_), .B(_1788_), .Y(_1800_) );
OAI21X1 OAI21X1_407 ( .A(_1799_), .B(_1788_), .C(_1800_), .Y(_1696_) );
INVX1 INVX1_266 ( .A(alu_inst_data_out_3_), .Y(_1801_) );
NAND2X1 NAND2X1_317 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_3_), .B(_1788_), .Y(_1802_) );
OAI21X1 OAI21X1_408 ( .A(_1801_), .B(_1788_), .C(_1802_), .Y(_1697_) );
INVX1 INVX1_267 ( .A(alu_inst_data_out_4_), .Y(_1803_) );
NAND2X1 NAND2X1_318 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_4_), .B(_1788_), .Y(_1804_) );
OAI21X1 OAI21X1_409 ( .A(_1803_), .B(_1788_), .C(_1804_), .Y(_1698_) );
INVX1 INVX1_268 ( .A(alu_inst_data_out_5_), .Y(_1805_) );
NAND2X1 NAND2X1_319 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_5_), .B(_1788_), .Y(_1806_) );
OAI21X1 OAI21X1_410 ( .A(_1805_), .B(_1788_), .C(_1806_), .Y(_1699_) );
INVX1 INVX1_269 ( .A(alu_inst_data_out_6_), .Y(_1807_) );
NAND2X1 NAND2X1_320 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_6_), .B(_1788_), .Y(_1808_) );
OAI21X1 OAI21X1_411 ( .A(_1807_), .B(_1788_), .C(_1808_), .Y(_1700_) );
INVX1 INVX1_270 ( .A(alu_inst_data_out_7_), .Y(_1809_) );
NAND2X1 NAND2X1_321 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_7_), .B(_1788_), .Y(_1810_) );
OAI21X1 OAI21X1_412 ( .A(_1809_), .B(_1788_), .C(_1810_), .Y(_1701_) );
INVX1 INVX1_271 ( .A(alu_inst_data_out_8_), .Y(_1811_) );
NAND2X1 NAND2X1_322 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_8_), .B(_1788_), .Y(_1812_) );
OAI21X1 OAI21X1_413 ( .A(_1811_), .B(_1788_), .C(_1812_), .Y(_1702_) );
INVX1 INVX1_272 ( .A(alu_inst_data_out_9_), .Y(_1813_) );
NAND2X1 NAND2X1_323 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_9_), .B(_1788_), .Y(_1814_) );
OAI21X1 OAI21X1_414 ( .A(_1813_), .B(_1788_), .C(_1814_), .Y(_1703_) );
INVX1 INVX1_273 ( .A(alu_inst_data_out_10_), .Y(_1815_) );
NAND2X1 NAND2X1_324 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_10_), .B(_1788_), .Y(_1816_) );
OAI21X1 OAI21X1_415 ( .A(_1815_), .B(_1788_), .C(_1816_), .Y(_1704_) );
INVX1 INVX1_274 ( .A(alu_inst_data_out_11_), .Y(_1817_) );
NAND2X1 NAND2X1_325 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_11_), .B(_1788_), .Y(_1818_) );
OAI21X1 OAI21X1_416 ( .A(_1817_), .B(_1788_), .C(_1818_), .Y(_1705_) );
INVX1 INVX1_275 ( .A(alu_inst_data_out_12_), .Y(_1819_) );
NAND2X1 NAND2X1_326 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_12_), .B(_1788_), .Y(_1820_) );
OAI21X1 OAI21X1_417 ( .A(_1819_), .B(_1788_), .C(_1820_), .Y(_1706_) );
INVX1 INVX1_276 ( .A(alu_inst_data_out_13_), .Y(_1821_) );
NAND2X1 NAND2X1_327 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_13_), .B(_1788_), .Y(_1822_) );
OAI21X1 OAI21X1_418 ( .A(_1821_), .B(_1788_), .C(_1822_), .Y(_1707_) );
INVX1 INVX1_277 ( .A(alu_inst_data_out_14_), .Y(_1823_) );
NAND2X1 NAND2X1_328 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_14_), .B(_1788_), .Y(_1824_) );
OAI21X1 OAI21X1_419 ( .A(_1823_), .B(_1788_), .C(_1824_), .Y(_1708_) );
INVX1 INVX1_278 ( .A(alu_inst_data_out_15_), .Y(_1825_) );
NAND2X1 NAND2X1_329 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_15_), .B(_1788_), .Y(_1826_) );
OAI21X1 OAI21X1_420 ( .A(_1825_), .B(_1788_), .C(_1826_), .Y(_1709_) );
INVX1 INVX1_279 ( .A(reg_file_inst_rd_data_out_0_), .Y(_1827_) );
NAND2X1 NAND2X1_330 ( .A(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_0_), .B(_1789_), .Y(_1828_) );
OAI21X1 OAI21X1_421 ( .A(_1827_), .B(_1789_), .C(_1828_), .Y(_1710_) );
INVX1 INVX1_280 ( .A(reg_file_inst_rd_data_out_1_), .Y(_1829_) );
NAND2X1 NAND2X1_331 ( .A(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_1_), .B(_1789_), .Y(_1830_) );
OAI21X1 OAI21X1_422 ( .A(_1829_), .B(_1789_), .C(_1830_), .Y(_1711_) );
INVX1 INVX1_281 ( .A(reg_file_inst_rd_data_out_2_), .Y(_1831_) );
NAND2X1 NAND2X1_332 ( .A(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_2_), .B(_1789_), .Y(_1832_) );
OAI21X1 OAI21X1_423 ( .A(_1831_), .B(_1789_), .C(_1832_), .Y(_1712_) );
INVX1 INVX1_282 ( .A(reg_file_inst_rd_data_out_3_), .Y(_1833_) );
NAND2X1 NAND2X1_333 ( .A(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_3_), .B(_1789_), .Y(_1834_) );
OAI21X1 OAI21X1_424 ( .A(_1833_), .B(_1789_), .C(_1834_), .Y(_1713_) );
INVX1 INVX1_283 ( .A(reg_file_inst_rd_data_out_4_), .Y(_1835_) );
NAND2X1 NAND2X1_334 ( .A(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_4_), .B(_1789_), .Y(_1836_) );
OAI21X1 OAI21X1_425 ( .A(_1835_), .B(_1789_), .C(_1836_), .Y(_1714_) );
INVX1 INVX1_284 ( .A(reg_file_inst_rd_data_out_5_), .Y(_1837_) );
NAND2X1 NAND2X1_335 ( .A(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_5_), .B(_1789_), .Y(_1838_) );
OAI21X1 OAI21X1_426 ( .A(_1837_), .B(_1789_), .C(_1838_), .Y(_1715_) );
INVX1 INVX1_285 ( .A(reg_file_inst_rd_data_out_6_), .Y(_1839_) );
NAND2X1 NAND2X1_336 ( .A(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_6_), .B(_1789_), .Y(_1840_) );
OAI21X1 OAI21X1_427 ( .A(_1839_), .B(_1789_), .C(_1840_), .Y(_1716_) );
INVX1 INVX1_286 ( .A(reg_file_inst_rd_data_out_7_), .Y(_1841_) );
NAND2X1 NAND2X1_337 ( .A(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_7_), .B(_1789_), .Y(_1842_) );
OAI21X1 OAI21X1_428 ( .A(_1841_), .B(_1789_), .C(_1842_), .Y(_1717_) );
DFFSR DFFSR_193 ( .CLK(ref_clk), .D(_1690_), .Q(sys_control_inst_sys_control_rx_inst_rf_addr_reg_0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_194 ( .CLK(ref_clk), .D(_1691_), .Q(sys_control_inst_sys_control_rx_inst_rf_addr_reg_1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_195 ( .CLK(ref_clk), .D(_1692_), .Q(sys_control_inst_sys_control_rx_inst_rf_addr_reg_2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_196 ( .CLK(ref_clk), .D(_1693_), .Q(sys_control_inst_sys_control_rx_inst_rf_addr_reg_3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_197 ( .CLK(ref_clk), .D(_1694_), .Q(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_198 ( .CLK(ref_clk), .D(_1695_), .Q(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_199 ( .CLK(ref_clk), .D(_1696_), .Q(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_200 ( .CLK(ref_clk), .D(_1697_), .Q(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_201 ( .CLK(ref_clk), .D(_1698_), .Q(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_202 ( .CLK(ref_clk), .D(_1699_), .Q(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_203 ( .CLK(ref_clk), .D(_1700_), .Q(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_204 ( .CLK(ref_clk), .D(_1701_), .Q(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_205 ( .CLK(ref_clk), .D(_1702_), .Q(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_8_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_206 ( .CLK(ref_clk), .D(_1703_), .Q(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_9_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_207 ( .CLK(ref_clk), .D(_1704_), .Q(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_10_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_208 ( .CLK(ref_clk), .D(_1705_), .Q(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_11_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_209 ( .CLK(ref_clk), .D(_1706_), .Q(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_12_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_210 ( .CLK(ref_clk), .D(_1707_), .Q(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_13_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_211 ( .CLK(ref_clk), .D(_1708_), .Q(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_14_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_212 ( .CLK(ref_clk), .D(_1709_), .Q(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_15_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_213 ( .CLK(ref_clk), .D(_1710_), .Q(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_214 ( .CLK(ref_clk), .D(_1711_), .Q(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_215 ( .CLK(ref_clk), .D(_1712_), .Q(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_216 ( .CLK(ref_clk), .D(_1713_), .Q(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_3_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_217 ( .CLK(ref_clk), .D(_1714_), .Q(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_4_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_218 ( .CLK(ref_clk), .D(_1715_), .Q(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_5_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_219 ( .CLK(ref_clk), .D(_1716_), .Q(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_6_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_220 ( .CLK(ref_clk), .D(_1717_), .Q(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_7_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_221 ( .CLK(ref_clk), .D(sys_control_inst_sys_control_rx_inst_next_state_0_), .Q(sys_control_inst_sys_control_rx_inst_current_state_0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_222 ( .CLK(ref_clk), .D(sys_control_inst_sys_control_rx_inst_next_state_1_), .Q(sys_control_inst_sys_control_rx_inst_current_state_1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_223 ( .CLK(ref_clk), .D(sys_control_inst_sys_control_rx_inst_next_state_2_), .Q(sys_control_inst_sys_control_rx_inst_current_state_2_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_224 ( .CLK(ref_clk), .D(sys_control_inst_sys_control_rx_inst_next_state_3_), .Q(sys_control_inst_sys_control_rx_inst_current_state_3_), .R(alu_inst_reset_n), .S(_true) );
INVX1 INVX1_287 ( .A(sys_control_inst_sys_control_tx_inst_current_state_1_), .Y(_1849_) );
INVX1 INVX1_288 ( .A(sys_control_inst_sys_control_tx_inst_current_state_2_), .Y(_1850_) );
NAND3X1 NAND3X1_215 ( .A(sys_control_inst_sys_control_tx_inst_current_state_0_), .B(_1849_), .C(_1850_), .Y(_1851_) );
INVX1 INVX1_289 ( .A(sys_control_inst_sys_control_tx_inst_current_state_0_), .Y(_1852_) );
NAND3X1 NAND3X1_216 ( .A(sys_control_inst_sys_control_tx_inst_current_state_2_), .B(_1849_), .C(_1852_), .Y(_1853_) );
NAND3X1 NAND3X1_217 ( .A(sys_control_inst_sys_control_tx_inst_current_state_1_), .B(_1852_), .C(_1850_), .Y(_1854_) );
NAND3X1 NAND3X1_218 ( .A(_1851_), .B(_1853_), .C(_1854_), .Y(data_synchronizer_inst_1_bus_enable_in) );
INVX1 INVX1_290 ( .A(_1854_), .Y(_1855_) );
NAND2X1 NAND2X1_338 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_0_), .B(_1855_), .Y(_1856_) );
INVX1 INVX1_291 ( .A(_1851_), .Y(_1857_) );
NAND2X1 NAND2X1_339 ( .A(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_0_), .B(_1857_), .Y(_1858_) );
INVX1 INVX1_292 ( .A(_1853_), .Y(_1859_) );
NAND2X1 NAND2X1_340 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_8_), .B(_1859_), .Y(_1860_) );
NAND3X1 NAND3X1_219 ( .A(_1856_), .B(_1858_), .C(_1860_), .Y(data_synchronizer_inst_1_unsync_data_in_0_) );
NAND2X1 NAND2X1_341 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_1_), .B(_1855_), .Y(_1861_) );
NAND2X1 NAND2X1_342 ( .A(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_1_), .B(_1857_), .Y(_1862_) );
NAND2X1 NAND2X1_343 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_9_), .B(_1859_), .Y(_1863_) );
NAND3X1 NAND3X1_220 ( .A(_1861_), .B(_1862_), .C(_1863_), .Y(data_synchronizer_inst_1_unsync_data_in_1_) );
NAND2X1 NAND2X1_344 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_2_), .B(_1855_), .Y(_1864_) );
NAND2X1 NAND2X1_345 ( .A(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_2_), .B(_1857_), .Y(_1865_) );
NAND2X1 NAND2X1_346 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_10_), .B(_1859_), .Y(_1866_) );
NAND3X1 NAND3X1_221 ( .A(_1864_), .B(_1865_), .C(_1866_), .Y(data_synchronizer_inst_1_unsync_data_in_2_) );
NAND2X1 NAND2X1_347 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_3_), .B(_1855_), .Y(_1867_) );
NAND2X1 NAND2X1_348 ( .A(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_3_), .B(_1857_), .Y(_1868_) );
NAND2X1 NAND2X1_349 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_11_), .B(_1859_), .Y(_1869_) );
NAND3X1 NAND3X1_222 ( .A(_1867_), .B(_1868_), .C(_1869_), .Y(data_synchronizer_inst_1_unsync_data_in_3_) );
NAND2X1 NAND2X1_350 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_4_), .B(_1855_), .Y(_1870_) );
NAND2X1 NAND2X1_351 ( .A(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_4_), .B(_1857_), .Y(_1871_) );
NAND2X1 NAND2X1_352 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_12_), .B(_1859_), .Y(_1872_) );
NAND3X1 NAND3X1_223 ( .A(_1870_), .B(_1871_), .C(_1872_), .Y(data_synchronizer_inst_1_unsync_data_in_4_) );
NAND2X1 NAND2X1_353 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_5_), .B(_1855_), .Y(_1873_) );
NAND2X1 NAND2X1_354 ( .A(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_5_), .B(_1857_), .Y(_1874_) );
NAND2X1 NAND2X1_355 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_13_), .B(_1859_), .Y(_1875_) );
NAND3X1 NAND3X1_224 ( .A(_1873_), .B(_1874_), .C(_1875_), .Y(data_synchronizer_inst_1_unsync_data_in_5_) );
NAND2X1 NAND2X1_356 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_6_), .B(_1855_), .Y(_1876_) );
NAND2X1 NAND2X1_357 ( .A(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_6_), .B(_1857_), .Y(_1877_) );
NAND2X1 NAND2X1_358 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_14_), .B(_1859_), .Y(_1878_) );
NAND3X1 NAND3X1_225 ( .A(_1876_), .B(_1877_), .C(_1878_), .Y(data_synchronizer_inst_1_unsync_data_in_6_) );
NAND2X1 NAND2X1_359 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_7_), .B(_1855_), .Y(_1879_) );
NAND2X1 NAND2X1_360 ( .A(sys_control_inst_sys_control_rx_inst_uart_rf_send_data_out_7_), .B(_1857_), .Y(_1880_) );
NAND2X1 NAND2X1_361 ( .A(sys_control_inst_sys_control_rx_inst_uart_alu_send_data_out_15_), .B(_1859_), .Y(_1881_) );
NAND3X1 NAND3X1_226 ( .A(_1879_), .B(_1880_), .C(_1881_), .Y(data_synchronizer_inst_1_unsync_data_in_7_) );
INVX1 INVX1_293 ( .A(bit_synchronizer_inst_sync_data_out), .Y(_1882_) );
NAND3X1 NAND3X1_227 ( .A(_1849_), .B(_1852_), .C(_1850_), .Y(_1883_) );
NOR2X1 NOR2X1_259 ( .A(sys_control_inst_sys_control_rx_inst_alu_data_store), .B(sys_control_inst_sys_control_rx_inst_rf_rd_store), .Y(_1884_) );
INVX1 INVX1_294 ( .A(_1884_), .Y(_1885_) );
NAND3X1 NAND3X1_228 ( .A(sys_control_inst_sys_control_tx_inst_current_state_1_), .B(sys_control_inst_sys_control_tx_inst_current_state_0_), .C(_1850_), .Y(_1886_) );
OAI22X1 OAI22X1_13 ( .A(_1882_), .B(_1886_), .C(_1883_), .D(_1885_), .Y(_1887_) );
AOI21X1 AOI21X1_139 ( .A(_1882_), .B(data_synchronizer_inst_1_bus_enable_in), .C(_1887_), .Y(_1888_) );
NAND2X1 NAND2X1_362 ( .A(_1882_), .B(data_synchronizer_inst_1_bus_enable_in), .Y(_1889_) );
NOR3X1 NOR3X1_21 ( .A(sys_control_inst_sys_control_tx_inst_current_state_1_), .B(sys_control_inst_sys_control_tx_inst_current_state_0_), .C(sys_control_inst_sys_control_tx_inst_current_state_2_), .Y(_1890_) );
NAND2X1 NAND2X1_363 ( .A(sys_control_inst_sys_control_tx_inst_current_state_1_), .B(sys_control_inst_sys_control_tx_inst_current_state_0_), .Y(_1891_) );
NOR2X1 NOR2X1_260 ( .A(sys_control_inst_sys_control_tx_inst_current_state_2_), .B(_1891_), .Y(_1892_) );
AOI22X1 AOI22X1_49 ( .A(_1890_), .B(_1884_), .C(_1892_), .D(bit_synchronizer_inst_sync_data_out), .Y(_1893_) );
INVX1 INVX1_295 ( .A(sys_control_inst_sys_control_rx_inst_rf_rd_store), .Y(_1894_) );
OAI21X1 OAI21X1_429 ( .A(_1894_), .B(_1883_), .C(_1854_), .Y(_1895_) );
NAND3X1 NAND3X1_229 ( .A(_1893_), .B(_1895_), .C(_1889_), .Y(_1896_) );
OAI21X1 OAI21X1_430 ( .A(_1852_), .B(_1888_), .C(_1896_), .Y(_1843_) );
OAI21X1 OAI21X1_431 ( .A(sys_control_inst_sys_control_rx_inst_rf_rd_store), .B(_1883_), .C(_1854_), .Y(_1846_) );
NAND3X1 NAND3X1_230 ( .A(_1893_), .B(_1846_), .C(_1889_), .Y(_1847_) );
OAI21X1 OAI21X1_432 ( .A(_1849_), .B(_1888_), .C(_1847_), .Y(_1844_) );
NAND3X1 NAND3X1_231 ( .A(_1892_), .B(_1893_), .C(_1889_), .Y(_1848_) );
OAI21X1 OAI21X1_433 ( .A(_1850_), .B(_1888_), .C(_1848_), .Y(_1845_) );
DFFSR DFFSR_225 ( .CLK(ref_clk), .D(_1843_), .Q(sys_control_inst_sys_control_tx_inst_current_state_0_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_226 ( .CLK(ref_clk), .D(_1844_), .Q(sys_control_inst_sys_control_tx_inst_current_state_1_), .R(alu_inst_reset_n), .S(_true) );
DFFSR DFFSR_227 ( .CLK(ref_clk), .D(_1845_), .Q(sys_control_inst_sys_control_tx_inst_current_state_2_), .R(alu_inst_reset_n), .S(_true) );
INVX1 INVX1_296 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_register_0_), .Y(_1900_) );
INVX1 INVX1_297 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_register_1_), .Y(_1901_) );
OAI21X1 OAI21X1_434 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_register_0_), .B(uart_top_inst_uart_rx_inst_data_sampling_inst_register_1_), .C(uart_top_inst_uart_rx_inst_data_sampling_inst_register_2_), .Y(_1902_) );
OAI21X1 OAI21X1_435 ( .A(_1900_), .B(_1901_), .C(_1902_), .Y(uart_top_inst_uart_rx_inst_data_sampling_inst_sampled_bit_out) );
INVX1 INVX1_298 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_2_), .Y(_1903_) );
NOR2X1 NOR2X1_261 ( .A(reg_file_inst_mem_2__5_), .B(_1903_), .Y(_1904_) );
NOR2X1 NOR2X1_262 ( .A(reg_file_inst_mem_2__3_), .B(reg_file_inst_mem_2__4_), .Y(_1905_) );
OR2X2 OR2X2_20 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_3_), .B(reg_file_inst_mem_2__6_), .Y(_1906_) );
NAND2X1 NAND2X1_364 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_3_), .B(reg_file_inst_mem_2__6_), .Y(_1907_) );
NAND2X1 NAND2X1_365 ( .A(_1907_), .B(_1906_), .Y(_1908_) );
AOI21X1 AOI21X1_140 ( .A(_1908_), .B(_1905_), .C(_1904_), .Y(_1909_) );
AOI22X1 AOI22X1_50 ( .A(_1903_), .B(reg_file_inst_mem_2__5_), .C(_1906_), .D(_1907_), .Y(_1910_) );
INVX1 INVX1_299 ( .A(_1910_), .Y(_1911_) );
NOR2X1 NOR2X1_263 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_1_), .B(reg_file_inst_mem_2__4_), .Y(_1912_) );
AND2X2 AND2X2_55 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_1_), .B(reg_file_inst_mem_2__4_), .Y(_1913_) );
OAI21X1 OAI21X1_436 ( .A(_1912_), .B(_1913_), .C(reg_file_inst_mem_2__3_), .Y(_1914_) );
INVX1 INVX1_300 ( .A(reg_file_inst_mem_2__3_), .Y(_1915_) );
OR2X2 OR2X2_21 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_1_), .B(reg_file_inst_mem_2__4_), .Y(_1916_) );
NAND2X1 NAND2X1_366 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_1_), .B(reg_file_inst_mem_2__4_), .Y(_1917_) );
NAND3X1 NAND3X1_232 ( .A(_1915_), .B(_1917_), .C(_1916_), .Y(_1918_) );
AND2X2 AND2X2_56 ( .A(_1918_), .B(_1914_), .Y(_1919_) );
AOI21X1 AOI21X1_141 ( .A(_1909_), .B(_1911_), .C(_1919_), .Y(_1920_) );
OR2X2 OR2X2_22 ( .A(reg_file_inst_mem_2__3_), .B(reg_file_inst_mem_2__4_), .Y(_1921_) );
XOR2X1 XOR2X1_48 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_3_), .B(reg_file_inst_mem_2__6_), .Y(_1922_) );
OAI22X1 OAI22X1_14 ( .A(_1903_), .B(reg_file_inst_mem_2__5_), .C(_1921_), .D(_1922_), .Y(_1923_) );
INVX1 INVX1_301 ( .A(reg_file_inst_mem_2__5_), .Y(_1924_) );
NOR2X1 NOR2X1_264 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_2_), .B(_1924_), .Y(_1925_) );
OAI21X1 OAI21X1_437 ( .A(_1925_), .B(_1922_), .C(_1905_), .Y(_1926_) );
XOR2X1 XOR2X1_49 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_0_), .B(reg_file_inst_mem_2__3_), .Y(_1927_) );
NOR2X1 NOR2X1_265 ( .A(reg_file_inst_mem_2__5_), .B(reg_file_inst_mem_2__6_), .Y(_1928_) );
INVX1 INVX1_302 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_4_), .Y(_1929_) );
NAND2X1 NAND2X1_367 ( .A(uart_top_inst_uart_rx_inst_counter_en), .B(_1929_), .Y(_1930_) );
AOI21X1 AOI21X1_142 ( .A(_1905_), .B(_1928_), .C(_1930_), .Y(_1931_) );
NAND2X1 NAND2X1_368 ( .A(_1927_), .B(_1931_), .Y(_1932_) );
AOI21X1 AOI21X1_143 ( .A(_1923_), .B(_1926_), .C(_1932_), .Y(_1933_) );
NAND3X1 NAND3X1_233 ( .A(rx_in), .B(_1933_), .C(_1920_), .Y(_1934_) );
NAND2X1 NAND2X1_369 ( .A(_1914_), .B(_1918_), .Y(_1935_) );
OAI21X1 OAI21X1_438 ( .A(_1910_), .B(_1923_), .C(_1935_), .Y(_1936_) );
AOI21X1 AOI21X1_144 ( .A(_1906_), .B(_1907_), .C(_1921_), .Y(_1937_) );
OAI22X1 OAI22X1_15 ( .A(_1921_), .B(_1910_), .C(_1904_), .D(_1937_), .Y(_1938_) );
XNOR2X1 XNOR2X1_23 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_0_), .B(reg_file_inst_mem_2__3_), .Y(_1939_) );
OR2X2 OR2X2_23 ( .A(reg_file_inst_mem_2__5_), .B(reg_file_inst_mem_2__6_), .Y(_1940_) );
INVX1 INVX1_303 ( .A(uart_top_inst_uart_rx_inst_counter_en), .Y(_1941_) );
NOR2X1 NOR2X1_266 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_4_), .B(_1941_), .Y(_1942_) );
OAI21X1 OAI21X1_439 ( .A(_1921_), .B(_1940_), .C(_1942_), .Y(_1943_) );
NOR2X1 NOR2X1_267 ( .A(_1939_), .B(_1943_), .Y(_1944_) );
NAND2X1 NAND2X1_370 ( .A(_1938_), .B(_1944_), .Y(_1945_) );
OAI21X1 OAI21X1_440 ( .A(_1936_), .B(_1945_), .C(uart_top_inst_uart_rx_inst_data_sampling_inst_register_0_), .Y(_1946_) );
NAND2X1 NAND2X1_371 ( .A(_1934_), .B(_1946_), .Y(_1897_) );
NOR2X1 NOR2X1_268 ( .A(_1930_), .B(_1927_), .Y(_1947_) );
AOI21X1 AOI21X1_145 ( .A(_1916_), .B(_1917_), .C(_1904_), .Y(_1948_) );
NAND3X1 NAND3X1_234 ( .A(_1910_), .B(_1948_), .C(_1947_), .Y(_1949_) );
NOR2X1 NOR2X1_269 ( .A(rx_in), .B(_1949_), .Y(_1950_) );
AOI21X1 AOI21X1_146 ( .A(_1901_), .B(_1949_), .C(_1950_), .Y(_1898_) );
XNOR2X1 XNOR2X1_24 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_2_), .B(reg_file_inst_mem_2__5_), .Y(_1951_) );
NAND2X1 NAND2X1_372 ( .A(reg_file_inst_mem_2__3_), .B(reg_file_inst_mem_2__4_), .Y(_1952_) );
INVX1 INVX1_304 ( .A(_1952_), .Y(_1953_) );
OAI22X1 OAI22X1_16 ( .A(_1951_), .B(_1953_), .C(_1925_), .D(_1908_), .Y(_1954_) );
NAND2X1 NAND2X1_373 ( .A(reg_file_inst_mem_2__5_), .B(reg_file_inst_mem_2__6_), .Y(_1955_) );
NOR2X1 NOR2X1_270 ( .A(_1952_), .B(_1955_), .Y(_1956_) );
NAND2X1 NAND2X1_374 ( .A(_1929_), .B(_1956_), .Y(_1957_) );
OAI21X1 OAI21X1_441 ( .A(_1903_), .B(reg_file_inst_mem_2__5_), .C(_1953_), .Y(_1958_) );
OAI21X1 OAI21X1_442 ( .A(_1958_), .B(_1922_), .C(_1957_), .Y(_1959_) );
NOR2X1 NOR2X1_271 ( .A(_1954_), .B(_1959_), .Y(_1960_) );
OAI21X1 OAI21X1_443 ( .A(_1952_), .B(_1955_), .C(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_4_), .Y(_1961_) );
NAND3X1 NAND3X1_235 ( .A(uart_top_inst_uart_rx_inst_counter_en), .B(_1961_), .C(_1927_), .Y(_1962_) );
NOR2X1 NOR2X1_272 ( .A(_1962_), .B(_1935_), .Y(_1963_) );
NAND3X1 NAND3X1_236 ( .A(rx_in), .B(_1963_), .C(_1960_), .Y(_1964_) );
OAI21X1 OAI21X1_444 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_2_), .B(_1924_), .C(_1922_), .Y(_1965_) );
OAI21X1 OAI21X1_445 ( .A(_1904_), .B(_1925_), .C(_1952_), .Y(_1966_) );
AOI21X1 AOI21X1_147 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_2_), .B(_1924_), .C(_1952_), .Y(_1967_) );
AOI22X1 AOI22X1_51 ( .A(_1929_), .B(_1956_), .C(_1908_), .D(_1967_), .Y(_1968_) );
NAND3X1 NAND3X1_237 ( .A(_1965_), .B(_1966_), .C(_1968_), .Y(_1969_) );
NOR2X1 NOR2X1_273 ( .A(_1941_), .B(_1939_), .Y(_1970_) );
NAND3X1 NAND3X1_238 ( .A(_1961_), .B(_1970_), .C(_1919_), .Y(_1971_) );
OAI21X1 OAI21X1_446 ( .A(_1969_), .B(_1971_), .C(uart_top_inst_uart_rx_inst_data_sampling_inst_register_2_), .Y(_1972_) );
NAND2X1 NAND2X1_375 ( .A(_1972_), .B(_1964_), .Y(_1899_) );
DFFSR DFFSR_228 ( .CLK(uart_clk), .D(_1897_), .Q(uart_top_inst_uart_rx_inst_data_sampling_inst_register_0_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_229 ( .CLK(uart_clk), .D(_1898_), .Q(uart_top_inst_uart_rx_inst_data_sampling_inst_register_1_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_230 ( .CLK(uart_clk), .D(_1899_), .Q(uart_top_inst_uart_rx_inst_data_sampling_inst_register_2_), .R(clk_divider_inst_reset_n), .S(_true) );
AND2X2 AND2X2_57 ( .A(data_synchronizer_inst_0_bus_enable_in), .B(uart_top_inst_uart_rx_inst_deserializer_inst_register_0_), .Y(data_synchronizer_inst_0_unsync_data_in_0_) );
AND2X2 AND2X2_58 ( .A(data_synchronizer_inst_0_bus_enable_in), .B(uart_top_inst_uart_rx_inst_deserializer_inst_register_1_), .Y(data_synchronizer_inst_0_unsync_data_in_1_) );
AND2X2 AND2X2_59 ( .A(data_synchronizer_inst_0_bus_enable_in), .B(uart_top_inst_uart_rx_inst_deserializer_inst_register_2_), .Y(data_synchronizer_inst_0_unsync_data_in_2_) );
AND2X2 AND2X2_60 ( .A(data_synchronizer_inst_0_bus_enable_in), .B(uart_top_inst_uart_rx_inst_deserializer_inst_register_3_), .Y(data_synchronizer_inst_0_unsync_data_in_3_) );
AND2X2 AND2X2_61 ( .A(data_synchronizer_inst_0_bus_enable_in), .B(uart_top_inst_uart_rx_inst_deserializer_inst_register_4_), .Y(data_synchronizer_inst_0_unsync_data_in_4_) );
AND2X2 AND2X2_62 ( .A(data_synchronizer_inst_0_bus_enable_in), .B(uart_top_inst_uart_rx_inst_deserializer_inst_register_5_), .Y(data_synchronizer_inst_0_unsync_data_in_5_) );
AND2X2 AND2X2_63 ( .A(data_synchronizer_inst_0_bus_enable_in), .B(uart_top_inst_uart_rx_inst_deserializer_inst_register_6_), .Y(data_synchronizer_inst_0_unsync_data_in_6_) );
AND2X2 AND2X2_64 ( .A(data_synchronizer_inst_0_bus_enable_in), .B(uart_top_inst_uart_rx_inst_deserializer_inst_register_7_), .Y(data_synchronizer_inst_0_unsync_data_in_7_) );
INVX1 INVX1_305 ( .A(uart_top_inst_uart_rx_inst_deserializer_inst_register_0_), .Y(_1981_) );
NAND2X1 NAND2X1_376 ( .A(uart_top_inst_uart_rx_inst_deserializer_inst_register_1_), .B(uart_top_inst_uart_rx_inst_deser_en), .Y(_1982_) );
OAI21X1 OAI21X1_447 ( .A(uart_top_inst_uart_rx_inst_deser_en), .B(_1981_), .C(_1982_), .Y(_1973_) );
INVX1 INVX1_306 ( .A(uart_top_inst_uart_rx_inst_deserializer_inst_register_1_), .Y(_1983_) );
NAND2X1 NAND2X1_377 ( .A(uart_top_inst_uart_rx_inst_deserializer_inst_register_2_), .B(uart_top_inst_uart_rx_inst_deser_en), .Y(_1984_) );
OAI21X1 OAI21X1_448 ( .A(uart_top_inst_uart_rx_inst_deser_en), .B(_1983_), .C(_1984_), .Y(_1974_) );
INVX1 INVX1_307 ( .A(uart_top_inst_uart_rx_inst_deserializer_inst_register_2_), .Y(_1985_) );
NAND2X1 NAND2X1_378 ( .A(uart_top_inst_uart_rx_inst_deserializer_inst_register_3_), .B(uart_top_inst_uart_rx_inst_deser_en), .Y(_1986_) );
OAI21X1 OAI21X1_449 ( .A(uart_top_inst_uart_rx_inst_deser_en), .B(_1985_), .C(_1986_), .Y(_1975_) );
INVX1 INVX1_308 ( .A(uart_top_inst_uart_rx_inst_deserializer_inst_register_3_), .Y(_1987_) );
NAND2X1 NAND2X1_379 ( .A(uart_top_inst_uart_rx_inst_deserializer_inst_register_4_), .B(uart_top_inst_uart_rx_inst_deser_en), .Y(_1988_) );
OAI21X1 OAI21X1_450 ( .A(uart_top_inst_uart_rx_inst_deser_en), .B(_1987_), .C(_1988_), .Y(_1976_) );
INVX1 INVX1_309 ( .A(uart_top_inst_uart_rx_inst_deserializer_inst_register_4_), .Y(_1989_) );
NAND2X1 NAND2X1_380 ( .A(uart_top_inst_uart_rx_inst_deserializer_inst_register_5_), .B(uart_top_inst_uart_rx_inst_deser_en), .Y(_1990_) );
OAI21X1 OAI21X1_451 ( .A(uart_top_inst_uart_rx_inst_deser_en), .B(_1989_), .C(_1990_), .Y(_1977_) );
INVX1 INVX1_310 ( .A(uart_top_inst_uart_rx_inst_deserializer_inst_register_5_), .Y(_1991_) );
NAND2X1 NAND2X1_381 ( .A(uart_top_inst_uart_rx_inst_deserializer_inst_register_6_), .B(uart_top_inst_uart_rx_inst_deser_en), .Y(_1992_) );
OAI21X1 OAI21X1_452 ( .A(uart_top_inst_uart_rx_inst_deser_en), .B(_1991_), .C(_1992_), .Y(_1978_) );
INVX1 INVX1_311 ( .A(uart_top_inst_uart_rx_inst_deserializer_inst_register_6_), .Y(_1993_) );
NAND2X1 NAND2X1_382 ( .A(uart_top_inst_uart_rx_inst_deserializer_inst_register_7_), .B(uart_top_inst_uart_rx_inst_deser_en), .Y(_1994_) );
OAI21X1 OAI21X1_453 ( .A(uart_top_inst_uart_rx_inst_deser_en), .B(_1993_), .C(_1994_), .Y(_1979_) );
INVX1 INVX1_312 ( .A(uart_top_inst_uart_rx_inst_deserializer_inst_register_7_), .Y(_1995_) );
NAND2X1 NAND2X1_383 ( .A(uart_top_inst_uart_rx_inst_deser_en), .B(uart_top_inst_uart_rx_inst_data_sampling_inst_sampled_bit_out), .Y(_1996_) );
OAI21X1 OAI21X1_454 ( .A(uart_top_inst_uart_rx_inst_deser_en), .B(_1995_), .C(_1996_), .Y(_1980_) );
DFFSR DFFSR_231 ( .CLK(uart_clk), .D(_1973_), .Q(uart_top_inst_uart_rx_inst_deserializer_inst_register_0_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_232 ( .CLK(uart_clk), .D(_1974_), .Q(uart_top_inst_uart_rx_inst_deserializer_inst_register_1_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_233 ( .CLK(uart_clk), .D(_1975_), .Q(uart_top_inst_uart_rx_inst_deserializer_inst_register_2_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_234 ( .CLK(uart_clk), .D(_1976_), .Q(uart_top_inst_uart_rx_inst_deserializer_inst_register_3_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_235 ( .CLK(uart_clk), .D(_1977_), .Q(uart_top_inst_uart_rx_inst_deserializer_inst_register_4_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_236 ( .CLK(uart_clk), .D(_1978_), .Q(uart_top_inst_uart_rx_inst_deserializer_inst_register_5_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_237 ( .CLK(uart_clk), .D(_1979_), .Q(uart_top_inst_uart_rx_inst_deserializer_inst_register_6_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_238 ( .CLK(uart_clk), .D(_1980_), .Q(uart_top_inst_uart_rx_inst_deserializer_inst_register_7_), .R(clk_divider_inst_reset_n), .S(_true) );
INVX1 INVX1_313 ( .A(uart_top_inst_uart_rx_inst_bit_count_0_), .Y(_2015_) );
INVX1 INVX1_314 ( .A(data_synchronizer_inst_0_bus_enable_in), .Y(_2016_) );
INVX1 INVX1_315 ( .A(uart_top_inst_uart_rx_inst_counter_en), .Y(_2017_) );
INVX1 INVX1_316 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_2_), .Y(_2018_) );
INVX1 INVX1_317 ( .A(reg_file_inst_mem_2__2_), .Y(_2019_) );
INVX1 INVX1_318 ( .A(reg_file_inst_mem_2__3_), .Y(_2020_) );
INVX1 INVX1_319 ( .A(reg_file_inst_mem_2__4_), .Y(_2021_) );
NAND3X1 NAND3X1_239 ( .A(_2019_), .B(_2020_), .C(_2021_), .Y(_2022_) );
OAI21X1 OAI21X1_455 ( .A(reg_file_inst_mem_2__2_), .B(reg_file_inst_mem_2__3_), .C(reg_file_inst_mem_2__4_), .Y(_2023_) );
NAND3X1 NAND3X1_240 ( .A(_2018_), .B(_2023_), .C(_2022_), .Y(_2024_) );
OAI21X1 OAI21X1_456 ( .A(reg_file_inst_mem_2__2_), .B(reg_file_inst_mem_2__3_), .C(_2021_), .Y(_2025_) );
NAND3X1 NAND3X1_241 ( .A(reg_file_inst_mem_2__4_), .B(_2019_), .C(_2020_), .Y(_2026_) );
NAND3X1 NAND3X1_242 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_2_), .B(_2025_), .C(_2026_), .Y(_2027_) );
NAND2X1 NAND2X1_384 ( .A(_2027_), .B(_2024_), .Y(_2028_) );
INVX1 INVX1_320 ( .A(reg_file_inst_mem_2__5_), .Y(_2029_) );
NAND2X1 NAND2X1_385 ( .A(_2029_), .B(_2022_), .Y(_2030_) );
NOR2X1 NOR2X1_274 ( .A(reg_file_inst_mem_2__2_), .B(reg_file_inst_mem_2__3_), .Y(_2031_) );
NAND3X1 NAND3X1_243 ( .A(_2021_), .B(reg_file_inst_mem_2__5_), .C(_2031_), .Y(_2032_) );
NAND3X1 NAND3X1_244 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_3_), .B(_2032_), .C(_2030_), .Y(_2033_) );
INVX1 INVX1_321 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_3_), .Y(_2034_) );
NOR2X1 NOR2X1_275 ( .A(reg_file_inst_mem_2__4_), .B(reg_file_inst_mem_2__5_), .Y(_2035_) );
NAND2X1 NAND2X1_386 ( .A(_2031_), .B(_2035_), .Y(_2036_) );
NAND2X1 NAND2X1_387 ( .A(reg_file_inst_mem_2__5_), .B(_2022_), .Y(_2037_) );
NAND3X1 NAND3X1_245 ( .A(_2034_), .B(_2036_), .C(_2037_), .Y(_2038_) );
NAND2X1 NAND2X1_388 ( .A(_2033_), .B(_2038_), .Y(_2039_) );
INVX1 INVX1_322 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_0_), .Y(_2040_) );
NAND2X1 NAND2X1_389 ( .A(reg_file_inst_mem_2__3_), .B(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_1_), .Y(_2041_) );
OR2X2 OR2X2_24 ( .A(reg_file_inst_mem_2__3_), .B(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_1_), .Y(_2042_) );
NAND3X1 NAND3X1_246 ( .A(_2040_), .B(_2041_), .C(_2042_), .Y(_2043_) );
AND2X2 AND2X2_65 ( .A(reg_file_inst_mem_2__3_), .B(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_1_), .Y(_2044_) );
NOR2X1 NOR2X1_276 ( .A(reg_file_inst_mem_2__3_), .B(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_1_), .Y(_2045_) );
OAI21X1 OAI21X1_457 ( .A(_2045_), .B(_2044_), .C(_2019_), .Y(_2046_) );
INVX1 INVX1_323 ( .A(reg_file_inst_mem_2__6_), .Y(_2047_) );
AOI22X1 AOI22X1_52 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_0_), .B(reg_file_inst_mem_2__2_), .C(_2047_), .D(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_4_), .Y(_2048_) );
NAND3X1 NAND3X1_247 ( .A(_2048_), .B(_2046_), .C(_2043_), .Y(_2049_) );
NOR2X1 NOR2X1_277 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_4_), .B(_2047_), .Y(_2050_) );
NAND3X1 NAND3X1_248 ( .A(_2031_), .B(_2035_), .C(_2050_), .Y(_2051_) );
OAI21X1 OAI21X1_458 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_4_), .B(_2047_), .C(_2036_), .Y(_2052_) );
AOI21X1 AOI21X1_148 ( .A(_2051_), .B(_2052_), .C(_2049_), .Y(_2053_) );
NAND3X1 NAND3X1_249 ( .A(_2028_), .B(_2039_), .C(_2053_), .Y(_2054_) );
OAI21X1 OAI21X1_459 ( .A(_2017_), .B(_2054_), .C(_2016_), .Y(_2055_) );
AND2X2 AND2X2_66 ( .A(_2046_), .B(_2048_), .Y(_2056_) );
NAND3X1 NAND3X1_250 ( .A(_2043_), .B(_2028_), .C(_2056_), .Y(_2057_) );
NAND3X1 NAND3X1_251 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_3_), .B(_2036_), .C(_2037_), .Y(_2058_) );
NAND3X1 NAND3X1_252 ( .A(_2034_), .B(_2032_), .C(_2030_), .Y(_2059_) );
NAND2X1 NAND2X1_390 ( .A(_2051_), .B(_2052_), .Y(_2060_) );
NAND3X1 NAND3X1_253 ( .A(_2058_), .B(_2059_), .C(_2060_), .Y(_2061_) );
NOR2X1 NOR2X1_278 ( .A(_2057_), .B(_2061_), .Y(_2062_) );
NOR2X1 NOR2X1_279 ( .A(data_synchronizer_inst_0_bus_enable_in), .B(_2017_), .Y(_2063_) );
NAND3X1 NAND3X1_254 ( .A(_2015_), .B(_2063_), .C(_2062_), .Y(_2064_) );
OAI21X1 OAI21X1_460 ( .A(_2015_), .B(_2055_), .C(_2064_), .Y(_1997_) );
INVX1 INVX1_324 ( .A(uart_top_inst_uart_rx_inst_bit_count_1_), .Y(_2065_) );
NAND2X1 NAND2X1_391 ( .A(_2016_), .B(_2017_), .Y(_2066_) );
OAI21X1 OAI21X1_461 ( .A(_2057_), .B(_2061_), .C(_2063_), .Y(_2067_) );
XNOR2X1 XNOR2X1_25 ( .A(uart_top_inst_uart_rx_inst_bit_count_0_), .B(uart_top_inst_uart_rx_inst_bit_count_1_), .Y(_2068_) );
NOR2X1 NOR2X1_280 ( .A(data_synchronizer_inst_0_bus_enable_in), .B(_2068_), .Y(_2069_) );
NAND3X1 NAND3X1_255 ( .A(_2066_), .B(_2069_), .C(_2067_), .Y(_2070_) );
OAI21X1 OAI21X1_462 ( .A(_2065_), .B(_2055_), .C(_2070_), .Y(_1998_) );
INVX1 INVX1_325 ( .A(uart_top_inst_uart_rx_inst_bit_count_2_), .Y(_2071_) );
NOR2X1 NOR2X1_281 ( .A(_2015_), .B(_2065_), .Y(_2072_) );
NAND2X1 NAND2X1_392 ( .A(uart_top_inst_uart_rx_inst_bit_count_2_), .B(_2072_), .Y(_2073_) );
INVX1 INVX1_326 ( .A(_2073_), .Y(_2074_) );
OAI21X1 OAI21X1_463 ( .A(uart_top_inst_uart_rx_inst_bit_count_2_), .B(_2072_), .C(_2016_), .Y(_2075_) );
NOR2X1 NOR2X1_282 ( .A(_2075_), .B(_2074_), .Y(_2076_) );
NAND3X1 NAND3X1_256 ( .A(_2066_), .B(_2076_), .C(_2067_), .Y(_2077_) );
OAI21X1 OAI21X1_464 ( .A(_2071_), .B(_2055_), .C(_2077_), .Y(_1999_) );
INVX1 INVX1_327 ( .A(uart_top_inst_uart_rx_inst_bit_count_3_), .Y(_2078_) );
NAND2X1 NAND2X1_393 ( .A(uart_top_inst_uart_rx_inst_bit_count_3_), .B(_2073_), .Y(_2079_) );
NAND2X1 NAND2X1_394 ( .A(_2078_), .B(_2074_), .Y(_2080_) );
AOI21X1 AOI21X1_149 ( .A(_2080_), .B(_2079_), .C(data_synchronizer_inst_0_bus_enable_in), .Y(_2081_) );
NAND3X1 NAND3X1_257 ( .A(_2066_), .B(_2081_), .C(_2067_), .Y(_2082_) );
OAI21X1 OAI21X1_465 ( .A(_2078_), .B(_2055_), .C(_2082_), .Y(_2000_) );
NAND3X1 NAND3X1_258 ( .A(_2016_), .B(_2040_), .C(_2054_), .Y(_2083_) );
MUX2X1 MUX2X1_3 ( .A(_2083_), .B(_2040_), .S(_2066_), .Y(_2001_) );
INVX1 INVX1_328 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_1_), .Y(_2006_) );
XNOR2X1 XNOR2X1_26 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_0_), .B(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_1_), .Y(_2007_) );
OAI22X1 OAI22X1_17 ( .A(_2006_), .B(_2066_), .C(_2007_), .D(_2067_), .Y(_2002_) );
NAND3X1 NAND3X1_259 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_0_), .B(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_1_), .C(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_2_), .Y(_2008_) );
OAI21X1 OAI21X1_466 ( .A(_2040_), .B(_2006_), .C(_2018_), .Y(_2009_) );
NAND2X1 NAND2X1_395 ( .A(_2008_), .B(_2009_), .Y(_2010_) );
OAI22X1 OAI22X1_18 ( .A(_2018_), .B(_2066_), .C(_2010_), .D(_2067_), .Y(_2003_) );
XOR2X1 XOR2X1_50 ( .A(_2008_), .B(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_3_), .Y(_2011_) );
OAI22X1 OAI22X1_19 ( .A(_2034_), .B(_2066_), .C(_2011_), .D(_2067_), .Y(_2004_) );
INVX1 INVX1_329 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_4_), .Y(_2012_) );
NOR2X1 NOR2X1_283 ( .A(_2034_), .B(_2008_), .Y(_2013_) );
XOR2X1 XOR2X1_51 ( .A(_2013_), .B(_2012_), .Y(_2014_) );
OAI22X1 OAI22X1_20 ( .A(_2012_), .B(_2066_), .C(_2014_), .D(_2067_), .Y(_2005_) );
DFFSR DFFSR_239 ( .CLK(uart_clk), .D(_1997_), .Q(uart_top_inst_uart_rx_inst_bit_count_0_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_240 ( .CLK(uart_clk), .D(_1998_), .Q(uart_top_inst_uart_rx_inst_bit_count_1_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_241 ( .CLK(uart_clk), .D(_1999_), .Q(uart_top_inst_uart_rx_inst_bit_count_2_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_242 ( .CLK(uart_clk), .D(_2000_), .Q(uart_top_inst_uart_rx_inst_bit_count_3_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_243 ( .CLK(uart_clk), .D(_2001_), .Q(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_0_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_244 ( .CLK(uart_clk), .D(_2002_), .Q(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_1_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_245 ( .CLK(uart_clk), .D(_2003_), .Q(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_2_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_246 ( .CLK(uart_clk), .D(_2004_), .Q(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_3_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_247 ( .CLK(uart_clk), .D(_2005_), .Q(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_4_), .R(clk_divider_inst_reset_n), .S(_true) );
INVX1 INVX1_330 ( .A(_false), .Y(_2084_) );
INVX1 INVX1_331 ( .A(uart_top_inst_uart_rx_inst_parity_check_inst_register), .Y(_2085_) );
NAND2X1 NAND2X1_396 ( .A(uart_top_inst_par_type_in), .B(_2085_), .Y(_2086_) );
INVX1 INVX1_332 ( .A(uart_top_inst_par_type_in), .Y(_2087_) );
NAND2X1 NAND2X1_397 ( .A(uart_top_inst_uart_rx_inst_parity_check_inst_register), .B(_2087_), .Y(_2088_) );
AOI21X1 AOI21X1_150 ( .A(_2086_), .B(_2088_), .C(_2084_), .Y(uart_top_inst_uart_rx_inst_par_err) );
DFFSR DFFSR_248 ( .CLK(uart_clk), .D(uart_top_inst_uart_rx_inst_data_sampling_inst_sampled_bit_out), .Q(uart_top_inst_uart_rx_inst_parity_check_inst_register), .R(clk_divider_inst_reset_n), .S(_true) );
INVX1 INVX1_333 ( .A(_false), .Y(_2089_) );
NOR2X1 NOR2X1_284 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_sampled_bit_out), .B(_2089_), .Y(uart_top_inst_uart_rx_inst_stop_check_inst_stp_err_out) );
AND2X2 AND2X2_67 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_sampled_bit_out), .B(uart_top_inst_uart_rx_inst_strt_check_inst_strt_chk_en_in), .Y(uart_top_inst_uart_rx_inst_strt_check_inst_strt_err_out) );
INVX1 INVX1_334 ( .A(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_0_), .Y(_2147_) );
NAND2X1 NAND2X1_398 ( .A(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_1_), .B(_2147_), .Y(_2148_) );
OAI21X1 OAI21X1_467 ( .A(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_2_), .B(_2147_), .C(_2148_), .Y(uart_top_inst_uart_rx_inst_counter_en) );
INVX1 INVX1_335 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_3_), .Y(_2149_) );
INVX1 INVX1_336 ( .A(reg_file_inst_mem_2__5_), .Y(_2150_) );
INVX1 INVX1_337 ( .A(reg_file_inst_mem_2__2_), .Y(_2151_) );
INVX1 INVX1_338 ( .A(reg_file_inst_mem_2__3_), .Y(_2152_) );
NAND2X1 NAND2X1_399 ( .A(_2151_), .B(_2152_), .Y(_2153_) );
OAI21X1 OAI21X1_468 ( .A(reg_file_inst_mem_2__4_), .B(_2153_), .C(_2150_), .Y(_2154_) );
INVX1 INVX1_339 ( .A(reg_file_inst_mem_2__4_), .Y(_2155_) );
NOR2X1 NOR2X1_285 ( .A(reg_file_inst_mem_2__2_), .B(reg_file_inst_mem_2__3_), .Y(_2156_) );
NAND3X1 NAND3X1_260 ( .A(_2155_), .B(reg_file_inst_mem_2__5_), .C(_2156_), .Y(_2157_) );
NAND3X1 NAND3X1_261 ( .A(_2149_), .B(_2157_), .C(_2154_), .Y(_2158_) );
NOR2X1 NOR2X1_286 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_1_), .B(reg_file_inst_mem_2__3_), .Y(_2159_) );
NAND2X1 NAND2X1_400 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_1_), .B(reg_file_inst_mem_2__3_), .Y(_2160_) );
INVX1 INVX1_340 ( .A(_2160_), .Y(_2161_) );
OAI21X1 OAI21X1_469 ( .A(_2159_), .B(_2161_), .C(_2151_), .Y(_2162_) );
INVX1 INVX1_341 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_0_), .Y(_2163_) );
INVX1 INVX1_342 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_1_), .Y(_2164_) );
NAND2X1 NAND2X1_401 ( .A(_2164_), .B(_2152_), .Y(_2165_) );
NAND3X1 NAND3X1_262 ( .A(_2163_), .B(_2160_), .C(_2165_), .Y(_2166_) );
AND2X2 AND2X2_68 ( .A(_2162_), .B(_2166_), .Y(_2167_) );
NAND2X1 NAND2X1_402 ( .A(_2155_), .B(_2150_), .Y(_2168_) );
INVX1 INVX1_343 ( .A(reg_file_inst_mem_2__6_), .Y(_2169_) );
NOR2X1 NOR2X1_287 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_4_), .B(_2169_), .Y(_2170_) );
OAI21X1 OAI21X1_470 ( .A(_2168_), .B(_2153_), .C(_2170_), .Y(_2171_) );
NAND3X1 NAND3X1_263 ( .A(_2171_), .B(_2158_), .C(_2167_), .Y(_2172_) );
AOI21X1 AOI21X1_151 ( .A(_2156_), .B(_2155_), .C(reg_file_inst_mem_2__5_), .Y(_2173_) );
INVX1 INVX1_344 ( .A(_2157_), .Y(_2174_) );
OAI21X1 OAI21X1_471 ( .A(_2173_), .B(_2174_), .C(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_3_), .Y(_2175_) );
OAI21X1 OAI21X1_472 ( .A(reg_file_inst_mem_2__2_), .B(reg_file_inst_mem_2__3_), .C(_2155_), .Y(_2176_) );
NAND3X1 NAND3X1_264 ( .A(reg_file_inst_mem_2__4_), .B(_2151_), .C(_2152_), .Y(_2177_) );
NAND2X1 NAND2X1_403 ( .A(_2176_), .B(_2177_), .Y(_2178_) );
NOR2X1 NOR2X1_288 ( .A(_2163_), .B(_2151_), .Y(_2179_) );
AOI21X1 AOI21X1_152 ( .A(_2178_), .B(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_2_), .C(_2179_), .Y(_2180_) );
INVX1 INVX1_345 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_2_), .Y(_2181_) );
INVX1 INVX1_346 ( .A(_2170_), .Y(_2182_) );
AND2X2 AND2X2_69 ( .A(_2177_), .B(_2176_), .Y(_2183_) );
INVX1 INVX1_347 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_4_), .Y(_2184_) );
OAI22X1 OAI22X1_21 ( .A(_2184_), .B(reg_file_inst_mem_2__6_), .C(_2168_), .D(_2153_), .Y(_2185_) );
AOI22X1 AOI22X1_53 ( .A(_2182_), .B(_2185_), .C(_2183_), .D(_2181_), .Y(_2186_) );
NAND3X1 NAND3X1_265 ( .A(_2180_), .B(_2175_), .C(_2186_), .Y(_2187_) );
NOR2X1 NOR2X1_289 ( .A(_2172_), .B(_2187_), .Y(_2188_) );
INVX1 INVX1_348 ( .A(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_2_), .Y(_2189_) );
NAND2X1 NAND2X1_404 ( .A(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_1_), .B(_2189_), .Y(_2190_) );
INVX1 INVX1_349 ( .A(uart_top_inst_uart_rx_inst_bit_count_1_), .Y(_2191_) );
INVX1 INVX1_350 ( .A(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_1_), .Y(_2192_) );
NAND2X1 NAND2X1_405 ( .A(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_0_), .B(_2189_), .Y(_2193_) );
NOR2X1 NOR2X1_290 ( .A(_2192_), .B(_2193_), .Y(_2194_) );
NOR2X1 NOR2X1_291 ( .A(uart_top_inst_uart_rx_inst_bit_count_0_), .B(uart_top_inst_uart_rx_inst_bit_count_2_), .Y(_2195_) );
AOI21X1 AOI21X1_153 ( .A(_2191_), .B(_2195_), .C(_2194_), .Y(_2196_) );
AOI21X1 AOI21X1_154 ( .A(_2196_), .B(uart_top_inst_uart_rx_inst_bit_count_3_), .C(_2190_), .Y(_2197_) );
AND2X2 AND2X2_70 ( .A(_2188_), .B(_2197_), .Y(uart_top_inst_uart_rx_inst_deser_en) );
NAND2X1 NAND2X1_406 ( .A(reg_file_inst_mem_2__4_), .B(reg_file_inst_mem_2__5_), .Y(_2198_) );
OR2X2 OR2X2_25 ( .A(_2198_), .B(_2169_), .Y(_2199_) );
OAI21X1 OAI21X1_473 ( .A(_2155_), .B(_2150_), .C(_2169_), .Y(_2200_) );
NAND2X1 NAND2X1_407 ( .A(_2200_), .B(_2199_), .Y(_2201_) );
NAND2X1 NAND2X1_408 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_3_), .B(_2201_), .Y(_2202_) );
AND2X2 AND2X2_71 ( .A(_2168_), .B(_2198_), .Y(_2203_) );
NAND2X1 NAND2X1_409 ( .A(_2164_), .B(_2155_), .Y(_2204_) );
NOR2X1 NOR2X1_292 ( .A(reg_file_inst_mem_2__3_), .B(_2163_), .Y(_2205_) );
NAND2X1 NAND2X1_410 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_1_), .B(reg_file_inst_mem_2__4_), .Y(_2206_) );
NAND2X1 NAND2X1_411 ( .A(_2206_), .B(_2204_), .Y(_2207_) );
OAI21X1 OAI21X1_474 ( .A(_2205_), .B(_2207_), .C(_2204_), .Y(_2208_) );
OAI21X1 OAI21X1_475 ( .A(_2203_), .B(_2208_), .C(_2181_), .Y(_2209_) );
NAND2X1 NAND2X1_412 ( .A(_2203_), .B(_2208_), .Y(_2210_) );
NAND2X1 NAND2X1_413 ( .A(_2210_), .B(_2209_), .Y(_2211_) );
NAND2X1 NAND2X1_414 ( .A(_2202_), .B(_2211_), .Y(_2212_) );
OAI21X1 OAI21X1_476 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_3_), .B(_2201_), .C(_2212_), .Y(_2213_) );
OAI21X1 OAI21X1_477 ( .A(_2169_), .B(_2198_), .C(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_4_), .Y(_2214_) );
NOR2X1 NOR2X1_293 ( .A(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_1_), .B(_2193_), .Y(_2093_) );
OAI21X1 OAI21X1_478 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_4_), .B(_2199_), .C(_2093_), .Y(_2094_) );
AOI21X1 AOI21X1_155 ( .A(_2213_), .B(_2214_), .C(_2094_), .Y(uart_top_inst_uart_rx_inst_strt_check_inst_strt_chk_en_in) );
OAI21X1 OAI21X1_479 ( .A(reg_file_inst_mem_2__3_), .B(reg_file_inst_mem_2__4_), .C(reg_file_inst_mem_2__5_), .Y(_2095_) );
INVX1 INVX1_351 ( .A(_2095_), .Y(_2096_) );
OAI21X1 OAI21X1_480 ( .A(_2149_), .B(_2096_), .C(_2184_), .Y(_2097_) );
OAI21X1 OAI21X1_481 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_3_), .B(_2095_), .C(_2182_), .Y(_2098_) );
NAND3X1 NAND3X1_266 ( .A(reg_file_inst_mem_2__6_), .B(_2097_), .C(_2098_), .Y(_2099_) );
OR2X2 OR2X2_26 ( .A(_2098_), .B(_2097_), .Y(_2100_) );
OAI21X1 OAI21X1_482 ( .A(reg_file_inst_mem_2__3_), .B(_2168_), .C(_2095_), .Y(_2101_) );
XOR2X1 XOR2X1_52 ( .A(_2101_), .B(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_2_), .Y(_2102_) );
INVX1 INVX1_352 ( .A(_2205_), .Y(_2103_) );
NAND3X1 NAND3X1_267 ( .A(_2163_), .B(reg_file_inst_mem_2__3_), .C(_2207_), .Y(_2104_) );
OAI21X1 OAI21X1_483 ( .A(_2103_), .B(_2207_), .C(_2104_), .Y(_2105_) );
INVX1 INVX1_353 ( .A(_2148_), .Y(_2106_) );
NAND2X1 NAND2X1_415 ( .A(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_2_), .B(_2106_), .Y(_2107_) );
OR2X2 OR2X2_27 ( .A(uart_top_inst_uart_rx_inst_stop_check_inst_stp_err_out), .B(uart_top_inst_uart_rx_inst_par_err), .Y(_2108_) );
NOR2X1 NOR2X1_294 ( .A(_2108_), .B(_2107_), .Y(_2109_) );
NAND3X1 NAND3X1_268 ( .A(_2105_), .B(_2109_), .C(_2102_), .Y(_2110_) );
AOI21X1 AOI21X1_156 ( .A(_2099_), .B(_2100_), .C(_2110_), .Y(data_synchronizer_inst_0_bus_enable_in) );
NOR2X1 NOR2X1_295 ( .A(_2173_), .B(_2174_), .Y(_2111_) );
NAND3X1 NAND3X1_269 ( .A(_2166_), .B(_2162_), .C(_2171_), .Y(_2112_) );
AOI21X1 AOI21X1_157 ( .A(_2111_), .B(_2149_), .C(_2112_), .Y(_2113_) );
AOI21X1 AOI21X1_158 ( .A(_2177_), .B(_2176_), .C(_2181_), .Y(_2114_) );
NAND3X1 NAND3X1_270 ( .A(_2181_), .B(_2176_), .C(_2177_), .Y(_2115_) );
NOR2X1 NOR2X1_296 ( .A(reg_file_inst_mem_2__4_), .B(reg_file_inst_mem_2__5_), .Y(_2116_) );
AOI22X1 AOI22X1_54 ( .A(uart_top_inst_uart_rx_inst_data_sampling_inst_edge_cnt_in_4_), .B(_2169_), .C(_2116_), .D(_2156_), .Y(_2117_) );
OAI21X1 OAI21X1_484 ( .A(_2170_), .B(_2117_), .C(_2115_), .Y(_2118_) );
NOR3X1 NOR3X1_22 ( .A(_2114_), .B(_2179_), .C(_2118_), .Y(_2119_) );
NAND3X1 NAND3X1_271 ( .A(_2175_), .B(_2119_), .C(_2113_), .Y(_2120_) );
INVX1 INVX1_354 ( .A(_2107_), .Y(_2121_) );
NOR2X1 NOR2X1_297 ( .A(uart_top_inst_uart_rx_inst_bit_count_3_), .B(uart_top_inst_uart_rx_inst_bit_count_2_), .Y(_2122_) );
NAND3X1 NAND3X1_272 ( .A(_2191_), .B(uart_top_inst_uart_rx_inst_bit_count_0_), .C(_2122_), .Y(_2123_) );
OAI21X1 OAI21X1_485 ( .A(uart_top_inst_uart_rx_inst_strt_check_inst_strt_err_out), .B(_2123_), .C(_2093_), .Y(_2124_) );
NAND2X1 NAND2X1_416 ( .A(uart_top_inst_uart_rx_inst_bit_count_0_), .B(_2191_), .Y(_2125_) );
INVX1 INVX1_355 ( .A(uart_top_inst_uart_rx_inst_bit_count_2_), .Y(_2126_) );
NAND2X1 NAND2X1_417 ( .A(uart_top_inst_uart_rx_inst_bit_count_3_), .B(_2126_), .Y(_2127_) );
OAI21X1 OAI21X1_486 ( .A(_2125_), .B(_2127_), .C(_2194_), .Y(_2128_) );
NOR2X1 NOR2X1_298 ( .A(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_2_), .B(_2148_), .Y(_2129_) );
NOR2X1 NOR2X1_299 ( .A(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_2_), .B(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_1_), .Y(_2130_) );
AND2X2 AND2X2_72 ( .A(_2130_), .B(_2147_), .Y(_2131_) );
NAND3X1 NAND3X1_273 ( .A(uart_top_inst_uart_rx_inst_bit_count_1_), .B(uart_top_inst_uart_rx_inst_bit_count_3_), .C(_2195_), .Y(_2132_) );
AOI22X1 AOI22X1_55 ( .A(_2131_), .B(rx_in), .C(_2129_), .D(_2132_), .Y(_2133_) );
NAND3X1 NAND3X1_274 ( .A(_2124_), .B(_2128_), .C(_2133_), .Y(_2134_) );
AOI21X1 AOI21X1_159 ( .A(_2120_), .B(_2121_), .C(_2134_), .Y(_2135_) );
OAI21X1 OAI21X1_487 ( .A(_2172_), .B(_2187_), .C(_2121_), .Y(_2136_) );
INVX1 INVX1_356 ( .A(_2134_), .Y(_2137_) );
AOI21X1 AOI21X1_160 ( .A(_2136_), .B(_2137_), .C(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_0_), .Y(_2138_) );
INVX1 INVX1_357 ( .A(uart_top_inst_par_en_in), .Y(_2139_) );
OAI21X1 OAI21X1_488 ( .A(_2147_), .B(_2139_), .C(_2130_), .Y(_2140_) );
NAND2X1 NAND2X1_418 ( .A(_2140_), .B(_2124_), .Y(_2141_) );
NOR2X1 NOR2X1_300 ( .A(rx_in), .B(_2107_), .Y(_2142_) );
AOI21X1 AOI21X1_161 ( .A(_2188_), .B(_2142_), .C(_2141_), .Y(_2143_) );
AOI21X1 AOI21X1_162 ( .A(_2143_), .B(_2135_), .C(_2138_), .Y(_2090_) );
NAND2X1 NAND2X1_419 ( .A(rx_in), .B(_2131_), .Y(_2144_) );
NAND2X1 NAND2X1_420 ( .A(_2144_), .B(_2124_), .Y(_2145_) );
OAI21X1 OAI21X1_489 ( .A(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_1_), .B(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_0_), .C(_2189_), .Y(_2146_) );
AOI21X1 AOI21X1_163 ( .A(_2135_), .B(_2146_), .C(_2145_), .Y(_2091_) );
OAI21X1 OAI21X1_490 ( .A(_2190_), .B(_2134_), .C(_2136_), .Y(_2092_) );
DFFSR DFFSR_249 ( .CLK(uart_clk), .D(_2090_), .Q(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_0_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_250 ( .CLK(uart_clk), .D(_2091_), .Q(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_1_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_251 ( .CLK(uart_clk), .D(_2092_), .Q(uart_top_inst_uart_rx_inst_uart_rx_fsm_inst_current_state_2_), .R(clk_divider_inst_reset_n), .S(_true) );
NAND3X1 NAND3X1_275 ( .A(uart_top_inst_uart_tx_inst_mux_inst_mux_sel_in_0_), .B(uart_top_inst_uart_tx_inst_mux_inst_mux_sel_in_1_), .C(uart_top_inst_uart_tx_inst_mux_inst_par_bit_in), .Y(_2215_) );
INVX1 INVX1_358 ( .A(uart_top_inst_uart_tx_inst_mux_inst_mux_sel_in_0_), .Y(_2216_) );
NAND3X1 NAND3X1_276 ( .A(uart_top_inst_uart_tx_inst_mux_inst_mux_sel_in_1_), .B(uart_top_inst_uart_tx_inst_mux_inst_data_in), .C(_2216_), .Y(_2217_) );
OR2X2 OR2X2_28 ( .A(uart_top_inst_uart_tx_inst_mux_inst_mux_sel_in_0_), .B(uart_top_inst_uart_tx_inst_mux_inst_mux_sel_in_1_), .Y(_2218_) );
NAND3X1 NAND3X1_277 ( .A(_2215_), .B(_2218_), .C(_2217_), .Y(_2313_) );
INVX1 INVX1_359 ( .A(data_synchronizer_inst_1_enable_pulse_out), .Y(_2220_) );
INVX1 INVX1_360 ( .A(uart_top_inst_uart_tx_inst_mux_inst_par_bit_in), .Y(_2221_) );
INVX1 INVX1_361 ( .A(data_synchronizer_inst_1_sync_data_out_5_), .Y(_2222_) );
INVX1 INVX1_362 ( .A(data_synchronizer_inst_1_sync_data_out_4_), .Y(_2223_) );
NAND2X1 NAND2X1_421 ( .A(_2222_), .B(_2223_), .Y(_2224_) );
NAND2X1 NAND2X1_422 ( .A(data_synchronizer_inst_1_sync_data_out_5_), .B(data_synchronizer_inst_1_sync_data_out_4_), .Y(_2225_) );
NAND2X1 NAND2X1_423 ( .A(data_synchronizer_inst_1_sync_data_out_3_), .B(data_synchronizer_inst_1_sync_data_out_2_), .Y(_2226_) );
OR2X2 OR2X2_29 ( .A(data_synchronizer_inst_1_sync_data_out_3_), .B(data_synchronizer_inst_1_sync_data_out_2_), .Y(_2227_) );
AOI22X1 AOI22X1_56 ( .A(_2227_), .B(_2226_), .C(_2224_), .D(_2225_), .Y(_2228_) );
NAND2X1 NAND2X1_424 ( .A(data_synchronizer_inst_1_sync_data_out_5_), .B(_2223_), .Y(_2229_) );
NAND2X1 NAND2X1_425 ( .A(data_synchronizer_inst_1_sync_data_out_4_), .B(_2222_), .Y(_2230_) );
XNOR2X1 XNOR2X1_27 ( .A(data_synchronizer_inst_1_sync_data_out_3_), .B(data_synchronizer_inst_1_sync_data_out_2_), .Y(_2231_) );
AOI21X1 AOI21X1_164 ( .A(_2229_), .B(_2230_), .C(_2231_), .Y(_2232_) );
NOR2X1 NOR2X1_301 ( .A(data_synchronizer_inst_1_sync_data_out_7_), .B(data_synchronizer_inst_1_sync_data_out_6_), .Y(_2233_) );
AND2X2 AND2X2_73 ( .A(data_synchronizer_inst_1_sync_data_out_7_), .B(data_synchronizer_inst_1_sync_data_out_6_), .Y(_2234_) );
OAI21X1 OAI21X1_491 ( .A(_2233_), .B(_2234_), .C(data_synchronizer_inst_1_sync_data_out_0_), .Y(_2235_) );
INVX1 INVX1_363 ( .A(data_synchronizer_inst_1_sync_data_out_0_), .Y(_2236_) );
OR2X2 OR2X2_30 ( .A(data_synchronizer_inst_1_sync_data_out_7_), .B(data_synchronizer_inst_1_sync_data_out_6_), .Y(_2237_) );
NAND2X1 NAND2X1_426 ( .A(data_synchronizer_inst_1_sync_data_out_7_), .B(data_synchronizer_inst_1_sync_data_out_6_), .Y(_2238_) );
NAND3X1 NAND3X1_278 ( .A(_2236_), .B(_2238_), .C(_2237_), .Y(_2239_) );
NAND2X1 NAND2X1_427 ( .A(_2235_), .B(_2239_), .Y(_2240_) );
OAI21X1 OAI21X1_492 ( .A(_2228_), .B(_2232_), .C(_2240_), .Y(_2241_) );
AOI21X1 AOI21X1_165 ( .A(_2224_), .B(_2225_), .C(_2231_), .Y(_2242_) );
AOI22X1 AOI22X1_57 ( .A(_2227_), .B(_2226_), .C(_2229_), .D(_2230_), .Y(_2243_) );
AND2X2 AND2X2_74 ( .A(_2239_), .B(_2235_), .Y(_2244_) );
OAI21X1 OAI21X1_493 ( .A(_2242_), .B(_2243_), .C(_2244_), .Y(_2245_) );
XNOR2X1 XNOR2X1_28 ( .A(uart_top_inst_par_type_in), .B(data_synchronizer_inst_1_sync_data_out_1_), .Y(_2246_) );
INVX1 INVX1_364 ( .A(_2246_), .Y(_2247_) );
NAND3X1 NAND3X1_279 ( .A(_2247_), .B(_2241_), .C(_2245_), .Y(_2248_) );
NAND2X1 NAND2X1_428 ( .A(_2241_), .B(_2245_), .Y(_2249_) );
AOI21X1 AOI21X1_166 ( .A(_2249_), .B(_2246_), .C(_2220_), .Y(_2250_) );
AOI22X1 AOI22X1_58 ( .A(_2220_), .B(_2221_), .C(_2250_), .D(_2248_), .Y(_2219_) );
DFFSR DFFSR_252 ( .CLK(clk_divider_inst_div_clk_out), .D(_2219_), .Q(uart_top_inst_uart_tx_inst_mux_inst_par_bit_in), .R(clk_divider_inst_reset_n), .S(_true) );
NAND3X1 NAND3X1_280 ( .A(uart_top_inst_uart_tx_inst_serializer_inst_counter_1_), .B(uart_top_inst_uart_tx_inst_serializer_inst_counter_0_), .C(uart_top_inst_uart_tx_inst_serializer_inst_counter_2_), .Y(_2262_) );
INVX1 INVX1_365 ( .A(_2262_), .Y(uart_top_inst_uart_tx_inst_ser_done) );
INVX1 INVX1_366 ( .A(uart_top_inst_uart_tx_inst_ser_en), .Y(_2263_) );
NAND3X1 NAND3X1_281 ( .A(_2263_), .B(uart_top_inst_uart_tx_inst_serializer_inst_counter_0_), .C(_2262_), .Y(_2264_) );
OAI21X1 OAI21X1_494 ( .A(_2263_), .B(uart_top_inst_uart_tx_inst_serializer_inst_counter_0_), .C(_2264_), .Y(_2251_) );
AOI21X1 AOI21X1_167 ( .A(uart_top_inst_uart_tx_inst_ser_en), .B(uart_top_inst_uart_tx_inst_serializer_inst_counter_0_), .C(uart_top_inst_uart_tx_inst_serializer_inst_counter_1_), .Y(_2265_) );
INVX1 INVX1_367 ( .A(uart_top_inst_uart_tx_inst_serializer_inst_counter_2_), .Y(_2266_) );
NAND2X1 NAND2X1_429 ( .A(uart_top_inst_uart_tx_inst_serializer_inst_counter_1_), .B(uart_top_inst_uart_tx_inst_serializer_inst_counter_0_), .Y(_2267_) );
AOI21X1 AOI21X1_168 ( .A(_2263_), .B(_2266_), .C(_2267_), .Y(_2268_) );
NOR2X1 NOR2X1_302 ( .A(_2265_), .B(_2268_), .Y(_2252_) );
OAI21X1 OAI21X1_495 ( .A(uart_top_inst_uart_tx_inst_ser_en), .B(uart_top_inst_uart_tx_inst_serializer_inst_counter_2_), .C(_2262_), .Y(_2269_) );
AOI21X1 AOI21X1_169 ( .A(_2266_), .B(_2267_), .C(_2269_), .Y(_2253_) );
INVX1 INVX1_368 ( .A(bit_synchronizer_inst_async_data_in), .Y(_2270_) );
NAND2X1 NAND2X1_430 ( .A(data_synchronizer_inst_1_enable_pulse_out), .B(_2270_), .Y(_2271_) );
NAND3X1 NAND3X1_282 ( .A(_2263_), .B(uart_top_inst_uart_tx_inst_mux_inst_data_in), .C(_2271_), .Y(_2272_) );
AOI22X1 AOI22X1_59 ( .A(uart_top_inst_uart_tx_inst_ser_en), .B(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_1_), .C(_2270_), .D(data_synchronizer_inst_1_enable_pulse_out), .Y(_2273_) );
INVX1 INVX1_369 ( .A(data_synchronizer_inst_1_enable_pulse_out), .Y(_2274_) );
NOR3X1 NOR3X1_23 ( .A(bit_synchronizer_inst_async_data_in), .B(data_synchronizer_inst_1_sync_data_out_0_), .C(_2274_), .Y(_2275_) );
OAI21X1 OAI21X1_496 ( .A(_2273_), .B(_2275_), .C(_2272_), .Y(_2254_) );
NAND3X1 NAND3X1_283 ( .A(_2263_), .B(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_1_), .C(_2271_), .Y(_2276_) );
AOI22X1 AOI22X1_60 ( .A(uart_top_inst_uart_tx_inst_ser_en), .B(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_2_), .C(_2270_), .D(data_synchronizer_inst_1_enable_pulse_out), .Y(_2277_) );
NOR3X1 NOR3X1_24 ( .A(bit_synchronizer_inst_async_data_in), .B(data_synchronizer_inst_1_sync_data_out_1_), .C(_2274_), .Y(_2278_) );
OAI21X1 OAI21X1_497 ( .A(_2277_), .B(_2278_), .C(_2276_), .Y(_2255_) );
NAND3X1 NAND3X1_284 ( .A(_2263_), .B(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_2_), .C(_2271_), .Y(_2279_) );
AOI22X1 AOI22X1_61 ( .A(uart_top_inst_uart_tx_inst_ser_en), .B(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_3_), .C(_2270_), .D(data_synchronizer_inst_1_enable_pulse_out), .Y(_2280_) );
NOR3X1 NOR3X1_25 ( .A(bit_synchronizer_inst_async_data_in), .B(data_synchronizer_inst_1_sync_data_out_2_), .C(_2274_), .Y(_2281_) );
OAI21X1 OAI21X1_498 ( .A(_2280_), .B(_2281_), .C(_2279_), .Y(_2256_) );
NAND3X1 NAND3X1_285 ( .A(_2263_), .B(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_3_), .C(_2271_), .Y(_2282_) );
AOI22X1 AOI22X1_62 ( .A(uart_top_inst_uart_tx_inst_ser_en), .B(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_4_), .C(_2270_), .D(data_synchronizer_inst_1_enable_pulse_out), .Y(_2283_) );
NOR3X1 NOR3X1_26 ( .A(bit_synchronizer_inst_async_data_in), .B(data_synchronizer_inst_1_sync_data_out_3_), .C(_2274_), .Y(_2284_) );
OAI21X1 OAI21X1_499 ( .A(_2283_), .B(_2284_), .C(_2282_), .Y(_2257_) );
NAND3X1 NAND3X1_286 ( .A(_2263_), .B(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_4_), .C(_2271_), .Y(_2285_) );
AOI22X1 AOI22X1_63 ( .A(uart_top_inst_uart_tx_inst_ser_en), .B(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_5_), .C(_2270_), .D(data_synchronizer_inst_1_enable_pulse_out), .Y(_2286_) );
NOR3X1 NOR3X1_27 ( .A(bit_synchronizer_inst_async_data_in), .B(data_synchronizer_inst_1_sync_data_out_4_), .C(_2274_), .Y(_2287_) );
OAI21X1 OAI21X1_500 ( .A(_2286_), .B(_2287_), .C(_2285_), .Y(_2258_) );
NAND3X1 NAND3X1_287 ( .A(_2263_), .B(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_5_), .C(_2271_), .Y(_2288_) );
AOI22X1 AOI22X1_64 ( .A(uart_top_inst_uart_tx_inst_ser_en), .B(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_6_), .C(_2270_), .D(data_synchronizer_inst_1_enable_pulse_out), .Y(_2289_) );
NOR3X1 NOR3X1_28 ( .A(bit_synchronizer_inst_async_data_in), .B(data_synchronizer_inst_1_sync_data_out_5_), .C(_2274_), .Y(_2290_) );
OAI21X1 OAI21X1_501 ( .A(_2289_), .B(_2290_), .C(_2288_), .Y(_2259_) );
NAND3X1 NAND3X1_288 ( .A(_2263_), .B(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_6_), .C(_2271_), .Y(_2291_) );
AOI22X1 AOI22X1_65 ( .A(uart_top_inst_uart_tx_inst_ser_en), .B(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_7_), .C(_2270_), .D(data_synchronizer_inst_1_enable_pulse_out), .Y(_2292_) );
NOR3X1 NOR3X1_29 ( .A(bit_synchronizer_inst_async_data_in), .B(data_synchronizer_inst_1_sync_data_out_6_), .C(_2274_), .Y(_2293_) );
OAI21X1 OAI21X1_502 ( .A(_2292_), .B(_2293_), .C(_2291_), .Y(_2260_) );
INVX1 INVX1_370 ( .A(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_7_), .Y(_2294_) );
INVX1 INVX1_371 ( .A(data_synchronizer_inst_1_sync_data_out_7_), .Y(_2295_) );
OAI21X1 OAI21X1_503 ( .A(bit_synchronizer_inst_async_data_in), .B(_2274_), .C(_2263_), .Y(_2296_) );
OAI22X1 OAI22X1_22 ( .A(_2295_), .B(_2271_), .C(_2294_), .D(_2296_), .Y(_2261_) );
DFFSR DFFSR_253 ( .CLK(clk_divider_inst_div_clk_out), .D(_2251_), .Q(uart_top_inst_uart_tx_inst_serializer_inst_counter_0_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_254 ( .CLK(clk_divider_inst_div_clk_out), .D(_2252_), .Q(uart_top_inst_uart_tx_inst_serializer_inst_counter_1_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_255 ( .CLK(clk_divider_inst_div_clk_out), .D(_2253_), .Q(uart_top_inst_uart_tx_inst_serializer_inst_counter_2_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_256 ( .CLK(clk_divider_inst_div_clk_out), .D(_2254_), .Q(uart_top_inst_uart_tx_inst_mux_inst_data_in), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_257 ( .CLK(clk_divider_inst_div_clk_out), .D(_2255_), .Q(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_1_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_258 ( .CLK(clk_divider_inst_div_clk_out), .D(_2256_), .Q(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_2_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_259 ( .CLK(clk_divider_inst_div_clk_out), .D(_2257_), .Q(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_3_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_260 ( .CLK(clk_divider_inst_div_clk_out), .D(_2258_), .Q(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_4_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_261 ( .CLK(clk_divider_inst_div_clk_out), .D(_2259_), .Q(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_5_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_262 ( .CLK(clk_divider_inst_div_clk_out), .D(_2260_), .Q(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_6_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_263 ( .CLK(clk_divider_inst_div_clk_out), .D(_2261_), .Q(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_7_), .R(clk_divider_inst_reset_n), .S(_true) );
INVX1 INVX1_372 ( .A(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_current_state_2_), .Y(_2298_) );
INVX1 INVX1_373 ( .A(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_current_state_0_), .Y(_2299_) );
NAND3X1 NAND3X1_289 ( .A(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_current_state_1_), .B(_2298_), .C(_2299_), .Y(_2300_) );
INVX1 INVX1_374 ( .A(_2300_), .Y(uart_top_inst_uart_tx_inst_ser_en) );
NAND2X1 NAND2X1_431 ( .A(uart_top_inst_uart_tx_inst_ser_done), .B(uart_top_inst_par_en_in), .Y(_2301_) );
INVX1 INVX1_375 ( .A(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_current_state_1_), .Y(_2302_) );
NAND3X1 NAND3X1_290 ( .A(data_synchronizer_inst_1_enable_pulse_out), .B(_2302_), .C(_2299_), .Y(_2303_) );
OAI21X1 OAI21X1_504 ( .A(_2301_), .B(_2300_), .C(_2303_), .Y(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_next_state_0_) );
NAND2X1 NAND2X1_432 ( .A(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_current_state_0_), .B(_2298_), .Y(_2304_) );
INVX1 INVX1_376 ( .A(uart_top_inst_uart_tx_inst_ser_done), .Y(_2305_) );
OAI21X1 OAI21X1_505 ( .A(_2305_), .B(uart_top_inst_par_en_in), .C(uart_top_inst_uart_tx_inst_ser_en), .Y(_2306_) );
OAI21X1 OAI21X1_506 ( .A(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_current_state_1_), .B(_2304_), .C(_2306_), .Y(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_next_state_1_) );
OR2X2 OR2X2_31 ( .A(_2305_), .B(uart_top_inst_par_en_in), .Y(_2307_) );
OAI22X1 OAI22X1_23 ( .A(_2302_), .B(_2304_), .C(_2300_), .D(_2307_), .Y(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_next_state_2_) );
INVX1 INVX1_377 ( .A(_2304_), .Y(uart_top_inst_uart_tx_inst_mux_inst_mux_sel_in_0_) );
NAND2X1 NAND2X1_433 ( .A(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_current_state_1_), .B(_2298_), .Y(_2308_) );
INVX1 INVX1_378 ( .A(_2308_), .Y(uart_top_inst_uart_tx_inst_mux_inst_mux_sel_in_1_) );
INVX1 INVX1_379 ( .A(_2303_), .Y(_2309_) );
OAI21X1 OAI21X1_507 ( .A(bit_synchronizer_inst_async_data_in), .B(_2309_), .C(_2298_), .Y(_2310_) );
NAND2X1 NAND2X1_434 ( .A(_2302_), .B(_2299_), .Y(_2311_) );
OAI21X1 OAI21X1_508 ( .A(_2311_), .B(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_next_state_0_), .C(bit_synchronizer_inst_async_data_in), .Y(_2312_) );
NAND2X1 NAND2X1_435 ( .A(_2310_), .B(_2312_), .Y(_2297_) );
DFFSR DFFSR_264 ( .CLK(clk_divider_inst_div_clk_out), .D(_2297_), .Q(bit_synchronizer_inst_async_data_in), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_265 ( .CLK(clk_divider_inst_div_clk_out), .D(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_next_state_0_), .Q(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_current_state_0_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_266 ( .CLK(clk_divider_inst_div_clk_out), .D(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_next_state_1_), .Q(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_current_state_1_), .R(clk_divider_inst_reset_n), .S(_true) );
DFFSR DFFSR_267 ( .CLK(clk_divider_inst_div_clk_out), .D(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_next_state_2_), .Q(uart_top_inst_uart_tx_inst_uart_tx_fsm_inst_current_state_2_), .R(clk_divider_inst_reset_n), .S(_true) );
BUFX2 BUFX2_1 ( .A(_2313_), .Y(tx_out) );
BUFX2 BUFX2_2 ( .A(uart_top_inst_par_en_in), .Y(reg_file_inst_mem_2__0_) );
BUFX2 BUFX2_3 ( .A(uart_top_inst_par_type_in), .Y(reg_file_inst_mem_2__1_) );
BUFX2 BUFX2_4 ( .A(clk_divider_inst_div_ratio_in_0_), .Y(reg_file_inst_mem_3__0_) );
BUFX2 BUFX2_5 ( .A(clk_divider_inst_div_ratio_in_1_), .Y(reg_file_inst_mem_3__1_) );
BUFX2 BUFX2_6 ( .A(clk_divider_inst_div_ratio_in_2_), .Y(reg_file_inst_mem_3__2_) );
BUFX2 BUFX2_7 ( .A(clk_divider_inst_div_ratio_in_3_), .Y(reg_file_inst_mem_3__3_) );
BUFX2 BUFX2_8 ( .A(clk_divider_inst_div_ratio_in_4_), .Y(reg_file_inst_mem_3__4_) );
BUFX2 BUFX2_9 ( .A(alu_inst_reset_n), .Y(reset_synchronizer_inst_0_ff_0_) );
BUFX2 BUFX2_10 ( .A(clk_divider_inst_reset_n), .Y(reset_synchronizer_inst_1_ff_0_) );
BUFX2 BUFX2_11 ( .A(uart_top_inst_uart_tx_inst_mux_inst_data_in), .Y(uart_top_inst_uart_tx_inst_serializer_inst_int_reg_0_) );
endmodule
