module \$_DLATCH_N_ (input CLK, input D, output Q);
  LATCH _TECHMAP_DLATCH_P (
    .D(D),
    .Q(Q),
    .CLK()
  );
endmodule